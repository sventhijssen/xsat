// Benchmark "top" written by ABC on Fri Mar 31 12:09:50 2023

module top ( 
    pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps, pd0, pe1,
    pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, px, ph1, pi0, pk2, py, ph2, pk1, pz, pi2, pj1, pk0, pl0, pm1,
    pn2, pl1, pm0, po2, pl2, pn0, po1, pm2, pn1, po0, pp0, pq1, pr2, pa,
    pp1, pq0, ps2, pb, pp2, pr0, ps1, pq2, pr1, ps0, pt0, pu1, pv2, pt1,
    pu0, pt2, pv0, pw1, pg, pu2, pv1, pw0, ph, px0, py1, pi, px1, py0, pz0,
    pk, pz1, pl, pm, pn, po,
    pc3, pd4, pe5, pb3, pd5, pe4, pa3, pf4, pg5, pf5, pg4, pa5, pg3, pa4,
    pf3, pb4, pc5, pe3, pb5, pc4, pd3, pk3, pl4, pm5, pj3, pl5, pm4, pi3,
    pn4, po5, ph3, pn5, po4, ph4, pi5, po3, ph5, pi4, pn3, pj4, pk5, pm3,
    pj5, pk4, pl3, ps3, pt4, pr3, pu4, pq3, pv4, pp3, pw4, pp4, pw3, pq4,
    pv3, pw2, pr4, pu3, ps4, pt3, pz2, pz3, px2, py3, px3, py2, px4, py4,
    pz4  );
  input  pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps,
    pd0, pe1, pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0,
    pw, ph0, pi1, pj2, px, ph1, pi0, pk2, py, ph2, pk1, pz, pi2, pj1, pk0,
    pl0, pm1, pn2, pl1, pm0, po2, pl2, pn0, po1, pm2, pn1, po0, pp0, pq1,
    pr2, pa, pp1, pq0, ps2, pb, pp2, pr0, ps1, pq2, pr1, ps0, pt0, pu1,
    pv2, pt1, pu0, pt2, pv0, pw1, pg, pu2, pv1, pw0, ph, px0, py1, pi, px1,
    py0, pz0, pk, pz1, pl, pm, pn, po;
  output pc3, pd4, pe5, pb3, pd5, pe4, pa3, pf4, pg5, pf5, pg4, pa5, pg3, pa4,
    pf3, pb4, pc5, pe3, pb5, pc4, pd3, pk3, pl4, pm5, pj3, pl5, pm4, pi3,
    pn4, po5, ph3, pn5, po4, ph4, pi5, po3, ph5, pi4, pn3, pj4, pk5, pm3,
    pj5, pk4, pl3, ps3, pt4, pr3, pu4, pq3, pv4, pp3, pw4, pp4, pw3, pq4,
    pv3, pw2, pr4, pu3, ps4, pt3, pz2, pz3, px2, py3, px3, py2, px4, py4,
    pz4;
  wire new_na1_, new_nb2_, new_np_, new_na0_, new_nc2_, new_nq_, new_nb0_,
    new_nc1_, new_nr_, new_na2_, new_nb1_, new_nc0_, new_ns_, new_nd0_,
    new_ne1_, new_nf2_, new_nt_, new_nd1_, new_ne0_, new_ng2_, new_nu_,
    new_nd2_, new_nf0_, new_ng1_, new_nv_, new_ne2_, new_nf1_, new_ng0_,
    new_nw_, new_nh0_, new_ni1_, new_nj2_, new_nx_, new_nh1_, new_ni0_,
    new_nk2_, new_ny_, new_nh2_, new_nk1_, new_nz_, new_ni2_, new_nj1_,
    new_nk0_, new_nl0_, new_nm1_, new_nn2_, new_nl1_, new_nm0_, new_no2_,
    new_nl2_, new_nn0_, new_no1_, new_nm2_, new_nn1_, new_no0_, new_np0_,
    new_nq1_, new_nr2_, new_na_, new_np1_, new_nq0_, new_ns2_, new_nb_,
    new_np2_, new_nr0_, new_ns1_, new_nq2_, new_nr1_, new_ns0_, new_nt0_,
    new_nu1_, new_nv2_, new_nt1_, new_nu0_, new_nt2_, new_nv0_, new_nw1_,
    new_ng_, new_nu2_, new_nv1_, new_nw0_, new_nh_, new_nx0_, new_ny1_,
    new_ni_, new_nx1_, new_ny0_, new_nz0_, new_nk_, new_nz1_, new_nl_,
    new_nm_, new_nn_, new_no_, new_ng3_, new_nr3_, new_n_n364_,
    new_n_n355_, new_n_n346_, new_n_n336_, new_n_n328_, new_nj4_,
    new_n_n312_, new_n_n304_, new_nu4_, new_n_n279_, new_n_n271_,
    new_n_n263_, new_n_n254_, new_n_n244_, new_n_n235_, new_n_n225_,
    new_n_n194_, new_n_n183_, new_n_n174_, new_n_n167_, new_n_n160_,
    new_nl9_, new_nv10_, new_nm13_, new_ny13_, new_nc14_, new_nh14_,
    new_n_n109_, new_n_n98_, new_nf3_, new_nh3_, new_ny3_, new_n_n356_,
    new_n_n345_, new_n_n337_, new_n_n327_, new_n_n321_, new_nm4_,
    new_n_n305_, new_n_n287_, new_n_n280_, new_n_n270_, new_nc5_,
    new_n_n253_, new_n_n245_, new_n_n234_, new_n_n226_, new_n_n203_,
    new_n_n182_, new_n_n175_, new_n_n166_, new_nx8_, new_nd10_, new_nu10_,
    new_np13_, new_n_n130_, new_n_n122_, new_ng14_, new_n_n108_,
    new_n_n99_, new_n_n369_, new_n_n363_, new_n_n353_, new_nb4_,
    new_n_n338_, new_ng4_, new_n_n319_, new_n_n314_, new_no4_, new_n_n286_,
    new_n_n278_, new_nz4_, new_n_n264_, new_n_n252_, new_ng5_, new_n_n237_,
    new_n_n227_, new_n_n202_, new_n_n192_, new_n_n176_, new_nm8_, new_nf9_,
    new_n_n154_, new_nn10_, new_nl11_, new_nl12_, new_nd14_, new_n_n116_,
    new_n_n111_, new_n_n100_, new_ne3_, new_n_n362_, new_n_n354_,
    new_n_n347_, new_n_n339_, new_n_n326_, new_n_n320_, new_n_n313_,
    new_n_n306_, new_n_n285_, new_nx4_, new_n_n272_, new_n_n265_,
    new_n_n251_, new_n_n243_, new_n_n236_, new_ni5_, new_n_n201_,
    new_n_n193_, new_n_n184_, new_no8_, new_n_n159_, new_n_n153_,
    new_nl10_, new_n_n136_, new_ni12_, new_n_n121_, new_nj14_, new_n_n110_,
    new_n_n101_, new_nk3_, new_nv3_, new_n_n340_, new_n_n325_, new_n_n301_,
    new_n_n293_, new_nf5_, new_n_n241_, new_n_n221_, new_n_n211_,
    new_n_n165_, new_n_n158_, new_n_n152_, new_nz10_, new_n_n142_,
    new_n_n120_, new_nk14_, new_n_n105_, new_n_n94_, new_n_n3_, new_nl3_,
    new_nu3_, new_n_n348_, new_n_n318_, new_n_n300_, new_ns4_, new_n_n250_,
    new_n_n242_, new_n_n220_, new_n_n212_, new_nw8_, new_ni9_, new_ny10_,
    new_na11_, new_n_n143_, new_ne14_, new_n_n115_, new_n_n104_,
    new_n_n95_, new_ni3_, new_nt3_, new_n_n357_, new_n_n311_, new_np4_,
    new_n_n294_, new_n_n233_, new_n_n223_, new_nj5_, new_n_n164_,
    new_ne10_, new_nx10_, new_nf14_, new_n_n114_, new_n_n107_, new_n_n96_,
    new_nj3_, new_ns3_, new_n_n365_, new_n_n303_, new_n_n302_, new_n_n295_,
    new_n_n232_, new_n_n224_, new_n_n222_, new_n_n157_, new_nf10_,
    new_n_n149_, new_n_n119_, new_nl14_, new_n_n106_, new_n_n97_, new_nc3_,
    new_no3_, new_nx3_, new_nz3_, new_n_n310_, new_n_n298_, new_n_n290_,
    new_nw4_, new_n_n273_, new_n_n217_, new_n_n207_, new_nk5_, new_n_n186_,
    new_nm5_, new_n_n147_, new_nk11_, new_nw11_, new_nd13_, new_nx13_,
    new_n_n124_, new_nb3_, new_np3_, new_nw3_, new_n_n349_, new_nk4_,
    new_n_n297_, new_nt4_, new_n_n281_, new_n_n274_, new_n_n216_,
    new_n_n208_, new_n_n196_, new_n_n187_, new_n_n169_, new_n_n146_,
    new_nj11_, new_nz11_, new_na13_, new_n_n131_, new_n_n125_, new_n_n0_,
    new_nm3_, new_n_n367_, new_n_n341_, new_n_n324_, new_nq4_, new_n_n291_,
    new_nb5_, new_ne5_, new_n_n219_, new_n_n209_, new_n_n195_, new_n_n178_,
    new_no5_, new_nc11_, new_ni11_, new_nc12_, new_nj13_, new_nw13_,
    new_n_n126_, new_n_n1_, new_nn3_, new_n_n368_, new_n_n332_,
    new_n_n331_, new_n_n299_, new_n_n292_, new_n_n266_, new_n_n259_,
    new_n_n218_, new_n_n210_, new_n_n185_, new_n_n177_, new_n_n170_,
    new_n_n148_, new_n_n141_, new_nf12_, new_ng13_, new_n_n132_, new_na14_,
    new_n_n2_, new_n_n370_, new_n_n361_, new_n_n352_, new_nc4_,
    new_n_n333_, new_ne4_, new_ni4_, new_n_n315_, new_n_n307_, new_nv4_,
    new_n_n276_, new_n_n268_, new_n_n260_, new_n_n258_, new_n_n248_,
    new_nh5_, new_n_n228_, new_n_n213_, new_n_n200_, new_n_n190_,
    new_n_n180_, new_n_n171_, new_n_n163_, new_n_n156_, new_n_n150_,
    new_nf11_, new_n_n137_, new_n_n135_, new_nr12_, new_n_n134_, new_nz13_,
    new_n_n113_, new_n_n102_, new_nx2_, new_nd3_, new_n_n360_, new_na4_,
    new_n_n342_, new_n_n334_, new_n_n330_, new_nh4_, new_nl4_, new_n_n308_,
    new_n_n284_, new_n_n277_, new_n_n267_, new_n_n261_, new_n_n257_,
    new_n_n249_, new_n_n238_, new_n_n229_, new_n_n204_, new_n_n199_,
    new_n_n191_, new_n_n179_, new_n_n172_, new_n_n168_, new_n_n155_,
    new_ng10_, new_n_n144_, new_n_n138_, new_nn11_, new_no12_, new_n_n133_,
    new_n_n127_, new_n_n112_, new_n_n103_, new_ny2_, new_n_n371_, new_nq3_,
    new_n_n359_, new_n_n350_, new_n_n344_, new_n_n335_, new_n_n329_,
    new_n_n322_, new_n_n317_, new_nn4_, new_nr4_, new_n_n288_, new_n_n283_,
    new_n_n275_, new_na5_, new_nd5_, new_n_n256_, new_n_n246_, new_n_n240_,
    new_n_n230_, new_n_n215_, new_n_n205_, new_n_n198_, new_n_n188_,
    new_n_n181_, new_n_n173_, new_nj8_, new_n_n161_, new_n_n151_,
    new_n_n145_, new_n_n139_, new_nq11_, new_nx12_, new_nu13_, new_n_n128_,
    new_nb14_, new_n_n117_, new_nz2_, new_n_n372_, new_n_n366_,
    new_n_n358_, new_n_n351_, new_n_n343_, new_nd4_, new_nf4_, new_n_n323_,
    new_n_n316_, new_n_n309_, new_n_n296_, new_n_n289_, new_n_n282_,
    new_ny4_, new_n_n269_, new_n_n262_, new_n_n255_, new_n_n247_,
    new_n_n239_, new_n_n231_, new_n_n214_, new_n_n206_, new_n_n197_,
    new_n_n189_, new_nl5_, new_nn5_, new_nk8_, new_n_n162_, new_nk9_,
    new_ne11_, new_n_n140_, new_nt11_, new_nu12_, new_nv13_, new_n_n129_,
    new_n_n123_, new_n_n118_, new_na3_, new_n_n88_, new_n_n77_, new_n_n66_,
    new_n_n55_, new_n_n44_, new_n_n89_, new_n_n76_, new_n_n67_, new_n_n54_,
    new_n_n45_, new_n_n90_, new_n_n75_, new_n_n64_, new_n_n57_, new_n_n46_,
    new_n_n91_, new_n_n74_, new_n_n65_, new_n_n56_, new_n_n47_, new_nw2_,
    new_n_n92_, new_n_n37_, new_n_n26_, new_n_n15_, new_n_n4_, new_n_n93_,
    new_n_n36_, new_n_n27_, new_n_n14_, new_n_n5_, new_n_n35_, new_n_n24_,
    new_n_n17_, new_n_n6_, new_n_n34_, new_n_n25_, new_n_n16_, new_n_n7_,
    new_n_n63_, new_n_n52_, new_n_n41_, new_n_n30_, new_n_n19_, new_n_n8_,
    new_n_n62_, new_n_n53_, new_n_n40_, new_n_n31_, new_n_n18_, new_n_n9_,
    new_n_n83_, new_n_n72_, new_n_n39_, new_n_n28_, new_n_n21_, new_n_n10_,
    new_n_n82_, new_n_n73_, new_n_n38_, new_n_n29_, new_n_n20_, new_n_n11_,
    new_n_n84_, new_n_n81_, new_n_n70_, new_n_n59_, new_n_n48_, new_n_n23_,
    new_n_n12_, new_n_n85_, new_n_n80_, new_n_n71_, new_n_n58_, new_n_n49_,
    new_n_n22_, new_n_n13_, new_n_n86_, new_n_n79_, new_n_n68_, new_n_n61_,
    new_n_n50_, new_n_n43_, new_n_n32_, new_n_n87_, new_n_n78_, new_n_n69_,
    new_n_n60_, new_n_n51_, new_n_n42_, new_n_n33_;
  assign new_na1_ = pa1;
  assign new_nb2_ = pb2;
  assign pc3 = new_nc3_;
  assign pd4 = new_nd4_;
  assign pe5 = new_ne5_;
  assign new_np_ = pp;
  assign new_na0_ = pa0;
  assign pb3 = new_nb3_;
  assign new_nc2_ = pc2;
  assign pd5 = new_nd5_;
  assign pe4 = new_ne4_;
  assign new_nq_ = pq;
  assign pa3 = new_na3_;
  assign new_nb0_ = pb0;
  assign new_nc1_ = pc1;
  assign pf4 = new_nf4_;
  assign pg5 = new_ng5_;
  assign new_nr_ = pr;
  assign new_na2_ = pa2;
  assign new_nb1_ = pb1;
  assign new_nc0_ = pc0;
  assign pf5 = new_nf5_;
  assign pg4 = new_ng4_;
  assign new_ns_ = ps;
  assign pa5 = new_na5_;
  assign new_nd0_ = pd0;
  assign new_ne1_ = pe1;
  assign new_nf2_ = pf2;
  assign pg3 = new_ng3_;
  assign new_nt_ = pt;
  assign pa4 = new_na4_;
  assign new_nd1_ = pd1;
  assign new_ne0_ = pe0;
  assign pf3 = new_nf3_;
  assign new_ng2_ = pg2;
  assign new_nu_ = pu;
  assign pb4 = new_nb4_;
  assign pc5 = new_nc5_;
  assign new_nd2_ = pd2;
  assign pe3 = new_ne3_;
  assign new_nf0_ = pf0;
  assign new_ng1_ = pg1;
  assign new_nv_ = pv;
  assign pb5 = new_nb5_;
  assign pc4 = new_nc4_;
  assign pd3 = new_nd3_;
  assign new_ne2_ = pe2;
  assign new_nf1_ = pf1;
  assign new_ng0_ = pg0;
  assign new_nw_ = pw;
  assign new_nh0_ = ph0;
  assign new_ni1_ = pi1;
  assign new_nj2_ = pj2;
  assign pk3 = new_nk3_;
  assign pl4 = new_nl4_;
  assign pm5 = new_nm5_;
  assign new_nx_ = px;
  assign new_nh1_ = ph1;
  assign new_ni0_ = pi0;
  assign pj3 = new_nj3_;
  assign new_nk2_ = pk2;
  assign pl5 = new_nl5_;
  assign pm4 = new_nm4_;
  assign new_ny_ = py;
  assign new_nh2_ = ph2;
  assign pi3 = new_ni3_;
  assign new_nk1_ = pk1;
  assign pn4 = new_nn4_;
  assign po5 = new_no5_;
  assign new_nz_ = pz;
  assign ph3 = new_nh3_;
  assign new_ni2_ = pi2;
  assign new_nj1_ = pj1;
  assign new_nk0_ = pk0;
  assign pn5 = new_nn5_;
  assign po4 = new_no4_;
  assign ph4 = new_nh4_;
  assign pi5 = new_ni5_;
  assign new_nl0_ = pl0;
  assign new_nm1_ = pm1;
  assign new_nn2_ = pn2;
  assign po3 = new_no3_;
  assign ph5 = new_nh5_;
  assign pi4 = new_ni4_;
  assign new_nl1_ = pl1;
  assign new_nm0_ = pm0;
  assign pn3 = new_nn3_;
  assign new_no2_ = po2;
  assign pj4 = new_nj4_;
  assign pk5 = new_nk5_;
  assign new_nl2_ = pl2;
  assign pm3 = new_nm3_;
  assign new_nn0_ = pn0;
  assign new_no1_ = po1;
  assign pj5 = new_nj5_;
  assign pk4 = new_nk4_;
  assign pl3 = new_nl3_;
  assign new_nm2_ = pm2;
  assign new_nn1_ = pn1;
  assign new_no0_ = po0;
  assign new_np0_ = pp0;
  assign new_nq1_ = pq1;
  assign new_nr2_ = pr2;
  assign ps3 = new_ns3_;
  assign pt4 = new_nt4_;
  assign new_na_ = pa;
  assign new_np1_ = pp1;
  assign new_nq0_ = pq0;
  assign pr3 = new_nr3_;
  assign new_ns2_ = ps2;
  assign pu4 = new_nu4_;
  assign new_nb_ = pb;
  assign new_np2_ = pp2;
  assign pq3 = new_nq3_;
  assign new_nr0_ = pr0;
  assign new_ns1_ = ps1;
  assign pv4 = new_nv4_;
  assign pp3 = new_np3_;
  assign new_nq2_ = pq2;
  assign new_nr1_ = pr1;
  assign new_ns0_ = ps0;
  assign pw4 = new_nw4_;
  assign pp4 = new_np4_;
  assign new_nt0_ = pt0;
  assign new_nu1_ = pu1;
  assign new_nv2_ = pv2;
  assign pw3 = new_nw3_;
  assign pq4 = new_nq4_;
  assign new_nt1_ = pt1;
  assign new_nu0_ = pu0;
  assign pv3 = new_nv3_;
  assign pw2 = new_nw2_;
  assign pr4 = new_nr4_;
  assign new_nt2_ = pt2;
  assign pu3 = new_nu3_;
  assign new_nv0_ = pv0;
  assign new_nw1_ = pw1;
  assign new_ng_ = pg;
  assign ps4 = new_ns4_;
  assign pt3 = new_nt3_;
  assign new_nu2_ = pu2;
  assign new_nv1_ = pv1;
  assign new_nw0_ = pw0;
  assign new_nh_ = ph;
  assign new_nx0_ = px0;
  assign new_ny1_ = py1;
  assign pz2 = new_nz2_;
  assign new_ni_ = pi;
  assign new_nx1_ = px1;
  assign new_ny0_ = py0;
  assign pz3 = new_nz3_;
  assign px2 = new_nx2_;
  assign py3 = new_ny3_;
  assign new_nz0_ = pz0;
  assign new_nk_ = pk;
  assign px3 = new_nx3_;
  assign py2 = new_ny2_;
  assign new_nz1_ = pz1;
  assign new_nl_ = pl;
  assign px4 = new_nx4_;
  assign new_nm_ = pm;
  assign py4 = new_ny4_;
  assign new_nn_ = pn;
  assign pz4 = new_nz4_;
  assign new_no_ = po;
  assign new_ng3_ = new_n_n58_ & new_n_n75_ & new_n_n5_;
  assign new_nr3_ = new_n_n75_ & new_nx0_;
  assign new_n_n364_ = new_n_n58_ & new_nl2_ & new_nm2_ & new_n_n104_;
  assign new_n_n355_ = new_np0_ & new_ng1_ & new_n_n58_;
  assign new_n_n346_ = new_n_n108_ & new_ni1_ & new_n_n58_;
  assign new_n_n336_ = new_n_n12_ & new_n_n11_ & new_n_n58_;
  assign new_n_n328_ = new_n_n62_ & new_nm1_;
  assign new_nj4_ = new_n_n320_ | new_n_n319_ | new_n_n318_;
  assign new_n_n312_ = new_n_n75_ & new_n_n40_ & new_n_n23_ & new_n_n80_;
  assign new_n_n304_ = new_ng0_ & new_n_n42_ & new_nq_ & new_n_n81_;
  assign new_nu4_ = new_n_n287_ | new_n_n286_ | new_n_n285_;
  assign new_n_n279_ = new_n_n75_ & new_n_n40_ & new_n_n34_ & new_n_n80_;
  assign new_n_n271_ = new_ng0_ & new_n_n42_ & new_nb0_ & new_n_n81_;
  assign new_n_n263_ = new_nj2_ & new_n_n75_ & new_n_n41_;
  assign new_n_n254_ = new_n_n103_ & new_n_n60_ & new_n_n44_;
  assign new_n_n244_ = new_nu2_ & new_n_n46_ & new_n_n45_;
  assign new_n_n235_ = new_n_n109_ & new_nd1_ & new_n_n48_;
  assign new_n_n225_ = new_n_n109_ & new_ne1_ & new_n_n49_;
  assign new_n_n194_ = new_nr2_ & new_n_n52_ & new_n_n58_;
  assign new_n_n183_ = new_ne1_ & new_n_n53_ & new_n_n58_ & new_n_n54_;
  assign new_n_n174_ = new_n_n58_ & new_ns2_ & new_n_n63_ & new_nl1_;
  assign new_n_n167_ = new_nt2_ & new_n_n79_;
  assign new_n_n160_ = new_n_n65_ & new_n_n67_;
  assign new_nl9_ = new_n_n68_ & new_n_n105_ & new_n_n112_;
  assign new_nv10_ = new_n_n149_ | new_ni0_;
  assign new_nm13_ = new_n_n108_ | new_n_n99_;
  assign new_ny13_ = new_n_n127_ | new_n_n129_ | new_n_n128_ | new_nc1_;
  assign new_nc14_ = new_n_n122_ | new_nc1_;
  assign new_nh14_ = new_n_n109_ | new_n_n112_ | new_n_n111_ | new_n_n105_;
  assign new_n_n109_ = ~new_nn2_;
  assign new_n_n98_ = ~new_nh2_;
  assign new_nf3_ = new_n_n368_ | new_n_n4_;
  assign new_nh3_ = new_n_n58_ & new_no0_ & new_n_n75_;
  assign new_ny3_ = new_n_n360_ | new_n_n359_ | new_n_n362_ | new_n_n361_ | new_n_n338_ | new_n_n358_ | new_n_n363_ | new_n_n336_;
  assign new_n_n356_ = new_n_n108_ & new_ng1_ & new_n_n58_;
  assign new_n_n345_ = new_nr0_ & new_ni1_ & new_n_n58_;
  assign new_n_n337_ = new_ns0_ & new_n_n11_ & new_n_n58_;
  assign new_n_n327_ = new_n_n62_ & new_n_n14_;
  assign new_n_n321_ = new_n_n75_ & new_n_n20_ & new_n_n40_ & new_n_n80_;
  assign new_nm4_ = new_n_n311_ | new_n_n310_ | new_n_n309_;
  assign new_n_n305_ = new_n_n75_ & new_n_n41_ & new_nv1_;
  assign new_n_n287_ = new_n_n75_ & new_n_n41_ & new_nb2_;
  assign new_n_n280_ = new_ng0_ & new_n_n42_ & new_ny_ & new_n_n81_;
  assign new_n_n270_ = new_n_n75_ & new_n_n40_ & new_n_n37_ & new_n_n80_;
  assign new_nc5_ = new_n_n262_ | new_n_n263_;
  assign new_n_n253_ = new_nl2_ & new_n_n46_ & new_n_n44_;
  assign new_n_n245_ = new_nm2_ & new_n_n46_ & new_n_n45_;
  assign new_n_n234_ = new_n_n111_ & new_nd1_ & new_n_n48_;
  assign new_n_n226_ = new_n_n111_ & new_np2_ & new_n_n49_;
  assign new_n_n203_ = new_n_n109_ & new_nd1_ & new_n_n51_;
  assign new_n_n182_ = new_nd1_ & new_n_n53_ & new_n_n58_ & new_n_n54_;
  assign new_n_n175_ = new_n_n58_ & new_n_n57_ & new_nt2_;
  assign new_n_n166_ = new_n_n63_ & new_nh0_;
  assign new_nx8_ = new_nc1_ | new_n_n160_ | new_n_n159_;
  assign new_nd10_ = new_n_n68_ | new_np2_ | new_no2_;
  assign new_nu10_ = new_n_n70_ | new_nh_ | new_ng_ | new_nk2_;
  assign new_np13_ = new_n_n108_ | new_n_n100_;
  assign new_n_n130_ = new_nm2_ & new_n_n104_;
  assign new_n_n122_ = new_n_n111_ & new_n_n109_;
  assign new_ng14_ = new_nr2_ & new_nq2_ & new_np2_;
  assign new_n_n108_ = ~new_ne1_;
  assign new_n_n99_ = ~new_ni2_;
  assign new_n_n369_ = new_nl0_ & new_n_n58_;
  assign new_n_n363_ = new_nn2_ & new_nf1_ & new_n_n58_;
  assign new_n_n353_ = new_np0_ & new_n_n11_ & new_n_n58_;
  assign new_nb4_ = new_n_n344_ | new_n_n359_ | new_n_n346_ | new_n_n345_ | new_n_n338_ | new_n_n343_ | new_n_n347_ | new_n_n336_;
  assign new_n_n338_ = new_n_n108_ & new_n_n11_ & new_n_n58_;
  assign new_ng4_ = new_n_n326_ | new_n_n325_ | new_n_n324_;
  assign new_n_n319_ = new_ng0_ & new_n_n42_ & new_nl_ & new_n_n81_;
  assign new_n_n314_ = new_n_n75_ & new_n_n41_ & new_ns1_;
  assign new_no4_ = new_n_n305_ | new_n_n304_ | new_n_n303_;
  assign new_n_n286_ = new_ng0_ & new_n_n42_ & new_nw_ & new_n_n81_;
  assign new_n_n278_ = new_n_n75_ & new_n_n41_ & new_ne2_;
  assign new_nz4_ = new_n_n272_ | new_n_n271_ | new_n_n270_;
  assign new_n_n264_ = new_n_n75_ & new_n_n40_ & new_n_n39_ & new_n_n80_;
  assign new_n_n252_ = new_nu2_ & new_n_n46_ & new_n_n44_;
  assign new_ng5_ = new_n_n239_ | new_n_n241_ | new_n_n240_ | new_n_n242_;
  assign new_n_n237_ = new_n_n109_ & new_ne1_ & new_n_n48_;
  assign new_n_n227_ = new_n_n109_ & new_np2_ & new_n_n49_;
  assign new_n_n202_ = new_n_n50_ & new_nd1_ & new_n_n51_;
  assign new_n_n192_ = new_n_n109_ & new_n_n53_ & new_n_n58_ & new_ne1_;
  assign new_n_n176_ = new_n_n58_ & new_n_n56_ & new_nt2_;
  assign new_nm8_ = new_n_n112_ & new_nr2_ & new_n_n64_;
  assign new_nf9_ = new_no2_ | new_nq2_ | new_np2_ | new_nr2_;
  assign new_n_n154_ = new_n_n66_ & new_n_n108_;
  assign new_nn10_ = new_n_n69_ | new_nn2_ | new_n_n108_ | new_n_n111_;
  assign new_nl11_ = new_n_n135_ | new_n_n136_;
  assign new_nl12_ = new_n_n108_ | new_n_n90_;
  assign new_nd14_ = new_nc1_ | new_n_n121_ | new_n_n120_;
  assign new_n_n116_ = new_n_n107_ & new_n_n106_;
  assign new_n_n111_ = ~new_no2_;
  assign new_n_n100_ = ~new_nj2_;
  assign new_ne3_ = new_n_n329_ | new_n_n369_;
  assign new_n_n362_ = new_n_n108_ & new_nf1_ & new_n_n58_;
  assign new_n_n354_ = new_n_n12_ & new_ng1_ & new_n_n58_;
  assign new_n_n347_ = new_nn2_ & new_ni1_ & new_n_n58_;
  assign new_n_n339_ = new_n_n12_ & new_nj1_ & new_n_n58_;
  assign new_n_n326_ = new_n_n75_ & new_nn1_ & new_n_n15_;
  assign new_n_n320_ = new_n_n75_ & new_n_n41_ & new_nq1_;
  assign new_n_n313_ = new_ng0_ & new_n_n42_ & new_nn_ & new_n_n81_;
  assign new_n_n306_ = new_n_n75_ & new_n_n40_ & new_n_n25_ & new_n_n80_;
  assign new_n_n285_ = new_n_n75_ & new_n_n40_ & new_n_n32_ & new_n_n80_;
  assign new_nx4_ = new_n_n278_ | new_n_n277_ | new_n_n276_;
  assign new_n_n272_ = new_n_n75_ & new_n_n41_ & new_ng2_;
  assign new_n_n265_ = new_ng0_ & new_n_n42_ & new_nd0_ & new_n_n81_;
  assign new_n_n251_ = new_n_n60_ & new_n_n46_ & new_n_n44_;
  assign new_n_n243_ = new_n_n60_ & new_n_n46_ & new_n_n45_;
  assign new_n_n236_ = new_n_n111_ & new_ne1_ & new_n_n48_;
  assign new_ni5_ = new_n_n224_ | new_n_n223_ | new_n_n226_ | new_n_n225_ | new_n_n214_ | new_n_n213_ | new_n_n227_ | new_n_n215_ | new_n_n221_ | new_n_n219_ | new_n_n222_ | new_n_n218_ | new_n_n220_ | new_n_n217_ | new_n_n216_;
  assign new_n_n201_ = new_n_n52_ & new_nd1_ & new_n_n51_;
  assign new_n_n193_ = new_nr2_ & new_n_n54_ & new_n_n58_;
  assign new_n_n184_ = new_n_n55_ & new_n_n53_ & new_n_n58_ & new_n_n52_;
  assign new_no8_ = new_n_n165_ | new_n_n108_ | new_no2_ | new_n_n109_;
  assign new_n_n159_ = new_n_n76_ & new_n_n65_;
  assign new_n_n153_ = new_n_n66_ & new_n_n69_;
  assign new_nl10_ = new_n_n68_ & new_n_n112_ & new_no2_ & new_n_n105_;
  assign new_n_n136_ = new_n_n80_ & new_ne1_;
  assign new_ni12_ = new_n_n108_ | new_n_n89_;
  assign new_n_n121_ = new_n_n112_ & new_n_n109_;
  assign new_nj14_ = new_ni0_ | new_n_n116_ | new_n_n115_;
  assign new_n_n110_ = ~new_nl14_;
  assign new_n_n101_ = ~new_nu0_;
  assign new_nk3_ = new_n_n58_ & new_nr0_ & new_n_n75_;
  assign new_nv3_ = new_n_n6_ | new_n_n368_ | new_n_n367_;
  assign new_n_n340_ = new_ns0_ & new_nj1_ & new_n_n58_;
  assign new_n_n325_ = new_n_n75_ & new_n_n17_ & new_n_n16_ & new_n_n80_;
  assign new_n_n301_ = new_ng0_ & new_n_n42_ & new_nr_ & new_n_n81_;
  assign new_n_n293_ = new_n_n75_ & new_n_n41_ & new_nz1_;
  assign new_nf5_ = new_n_n247_ | new_n_n246_ | new_n_n249_ | new_n_n248_ | new_n_n245_ | new_n_n244_ | new_n_n250_ | new_n_n243_;
  assign new_n_n241_ = new_n_n47_ & new_ne1_;
  assign new_n_n221_ = new_n_n111_ & new_nd1_ & new_n_n49_;
  assign new_n_n211_ = new_n_n109_ & new_nq2_ & new_n_n51_;
  assign new_n_n165_ = new_n_n105_ & new_n_n73_;
  assign new_n_n158_ = new_n_n80_ & new_n_n75_;
  assign new_n_n152_ = new_n_n75_ & new_n_n67_;
  assign new_nz10_ = new_n_n140_ | new_n_n139_ | new_n_n137_;
  assign new_n_n142_ = new_n_n75_ & new_n_n74_ & new_np1_;
  assign new_n_n120_ = new_n_n112_ & new_n_n111_;
  assign new_nk14_ = new_n_n108_ | new_n_n109_ | new_n_n110_;
  assign new_n_n105_ = ~new_nq2_;
  assign new_n_n94_ = ~new_nd2_;
  assign new_n_n3_ = ~new_nx8_;
  assign new_nl3_ = new_n_n58_ & new_ns0_ & new_n_n75_;
  assign new_nu3_ = new_n_n75_ & new_na1_;
  assign new_n_n348_ = new_nq0_ & new_n_n11_ & new_n_n58_;
  assign new_n_n318_ = new_n_n75_ & new_n_n40_ & new_n_n21_ & new_n_n80_;
  assign new_n_n300_ = new_n_n75_ & new_n_n40_ & new_n_n27_ & new_n_n80_;
  assign new_ns4_ = new_n_n293_ | new_n_n292_ | new_n_n291_;
  assign new_n_n250_ = new_n_n103_ & new_nm2_ & new_n_n45_;
  assign new_n_n242_ = new_n_n47_ & new_nn2_;
  assign new_n_n220_ = new_n_n112_ & new_nd1_ & new_n_n49_;
  assign new_n_n212_ = new_n_n111_ & new_nq2_ & new_n_n51_;
  assign new_nw8_ = new_n_n161_ | new_n_n163_ | new_n_n162_ | new_n_n164_;
  assign new_ni9_ = new_n_n157_ | new_n_n158_;
  assign new_ny10_ = new_n_n108_ | new_no1_;
  assign new_na11_ = new_n_n77_ | new_n_n76_;
  assign new_n_n143_ = new_n_n75_ & new_n_n108_ & new_n_n74_;
  assign new_ne14_ = new_np2_ & new_nq2_;
  assign new_n_n115_ = new_nu0_ & new_n_n107_;
  assign new_n_n104_ = ~new_nk2_;
  assign new_n_n95_ = ~new_ne2_;
  assign new_ni3_ = new_n_n58_ & new_np0_ & new_n_n75_;
  assign new_nt3_ = new_n_n75_ & new_nz0_;
  assign new_n_n357_ = new_nn2_ & new_ng1_ & new_n_n58_;
  assign new_n_n311_ = new_n_n75_ & new_n_n41_ & new_nt1_;
  assign new_np4_ = new_n_n302_ | new_n_n301_ | new_n_n300_;
  assign new_n_n294_ = new_n_n75_ & new_n_n40_ & new_n_n29_ & new_n_n80_;
  assign new_n_n233_ = new_n_n109_ & new_n_n55_ & new_n_n48_;
  assign new_n_n223_ = new_n_n112_ & new_ne1_ & new_n_n49_;
  assign new_nj5_ = new_n_n209_ | new_n_n208_ | new_n_n211_ | new_n_n210_ | new_n_n199_ | new_n_n198_ | new_n_n212_ | new_n_n200_ | new_n_n201_ | new_n_n203_ | new_n_n197_ | new_n_n202_ | new_n_n205_ | new_n_n204_ | new_n_n207_ | new_n_n206_;
  assign new_n_n164_ = new_nm1_ & new_ng_;
  assign new_ne10_ = new_n_n73_ & new_n_n105_;
  assign new_nx10_ = new_nl2_ & new_nm2_;
  assign new_nf14_ = new_n_n117_ | new_n_n119_ | new_n_n118_ | new_nc1_;
  assign new_n_n114_ = new_ni_ & new_n_n111_ & new_nr2_ & new_n_n112_;
  assign new_n_n107_ = ~new_nu2_;
  assign new_n_n96_ = ~new_nf2_;
  assign new_nj3_ = new_n_n58_ & new_nq0_ & new_n_n75_;
  assign new_ns3_ = new_n_n75_ & new_ny0_;
  assign new_n_n365_ = new_nd1_ & new_n_n58_;
  assign new_n_n303_ = new_n_n75_ & new_n_n40_ & new_n_n26_ & new_n_n80_;
  assign new_n_n302_ = new_n_n75_ & new_n_n41_ & new_nw1_;
  assign new_n_n295_ = new_ng0_ & new_n_n42_ & new_nt_ & new_n_n81_;
  assign new_n_n232_ = new_n_n111_ & new_n_n55_ & new_n_n48_;
  assign new_n_n224_ = new_n_n111_ & new_ne1_ & new_n_n49_;
  assign new_n_n222_ = new_n_n109_ & new_nd1_ & new_n_n49_;
  assign new_n_n157_ = new_n_n75_ & new_nv2_ & new_ng0_;
  assign new_nf10_ = new_n_n151_ | new_n_n152_;
  assign new_n_n149_ = new_ng0_ & new_nv2_;
  assign new_n_n119_ = new_n_n105_ & new_n_n109_;
  assign new_nl14_ = new_n_n113_ | new_n_n114_;
  assign new_n_n106_ = ~new_nb_;
  assign new_n_n97_ = ~new_ng2_;
  assign new_nc3_ = new_n_n371_ | new_n_n372_;
  assign new_no3_ = new_na_ & new_n_n75_;
  assign new_nx3_ = new_n_n366_ | new_n_n365_ | new_n_n364_;
  assign new_nz3_ = new_n_n354_ | new_n_n359_ | new_n_n356_ | new_n_n355_ | new_n_n338_ | new_n_n353_ | new_n_n357_ | new_n_n336_;
  assign new_n_n310_ = new_ng0_ & new_n_n42_ & new_no_ & new_n_n81_;
  assign new_n_n298_ = new_ng0_ & new_n_n42_ & new_ns_ & new_n_n81_;
  assign new_n_n290_ = new_n_n75_ & new_n_n41_ & new_na2_;
  assign new_nw4_ = new_n_n281_ | new_n_n280_ | new_n_n279_;
  assign new_n_n273_ = new_n_n75_ & new_n_n40_ & new_n_n36_ & new_n_n80_;
  assign new_n_n217_ = new_n_n112_ & new_n_n55_ & new_n_n49_;
  assign new_n_n207_ = new_n_n109_ & new_ne1_ & new_n_n51_;
  assign new_nk5_ = new_n_n193_ | new_n_n192_ | new_n_n195_ | new_n_n194_ | new_n_n183_ | new_n_n182_ | new_n_n196_ | new_n_n184_ | new_n_n185_ | new_n_n187_ | new_n_n181_ | new_n_n186_ | new_n_n189_ | new_n_n188_ | new_n_n191_ | new_n_n190_;
  assign new_n_n186_ = new_ne1_ & new_n_n53_ & new_n_n58_ & new_n_n52_;
  assign new_nm5_ = new_n_n176_ | new_n_n175_ | new_n_n174_;
  assign new_n_n147_ = new_n_n79_ & new_ng0_ & new_nm1_ & new_nv2_;
  assign new_nk11_ = new_n_n137_ | new_n_n139_ | new_n_n138_ | new_n_n140_;
  assign new_nw11_ = new_n_n108_ | new_n_n85_;
  assign new_nd13_ = new_n_n108_ | new_n_n96_;
  assign new_nx13_ = new_nc1_ | new_n_n131_ | new_n_n130_;
  assign new_n_n124_ = new_n_n104_ & new_nl2_ & new_nm2_ & new_nn2_;
  assign new_nb3_ = ~new_nk1_;
  assign new_np3_ = new_n_n75_ & new_nv0_;
  assign new_nw3_ = new_n_n10_ & new_nv2_;
  assign new_n_n349_ = new_n_n12_ & new_nh1_ & new_n_n58_;
  assign new_nk4_ = new_n_n317_ | new_n_n316_ | new_n_n315_;
  assign new_n_n297_ = new_n_n75_ & new_n_n40_ & new_n_n28_ & new_n_n80_;
  assign new_nt4_ = new_n_n290_ | new_n_n289_ | new_n_n288_;
  assign new_n_n281_ = new_n_n75_ & new_n_n41_ & new_nd2_;
  assign new_n_n274_ = new_ng0_ & new_n_n42_ & new_na0_ & new_n_n81_;
  assign new_n_n216_ = new_np2_ & new_n_n52_ & new_n_n49_;
  assign new_n_n208_ = new_n_n111_ & new_ne1_ & new_n_n51_;
  assign new_n_n196_ = new_n_n109_ & new_nr2_ & new_n_n58_;
  assign new_n_n187_ = new_n_n111_ & new_n_n53_ & new_n_n58_ & new_n_n55_;
  assign new_n_n169_ = new_n_n61_ & new_n_n62_;
  assign new_n_n146_ = new_nv2_ & new_ng_ & new_nm1_ & new_ng0_;
  assign new_nj11_ = new_n_n108_ | new_n_n78_;
  assign new_nz11_ = new_n_n108_ | new_n_n86_;
  assign new_na13_ = new_n_n108_ | new_n_n95_;
  assign new_n_n131_ = new_n_n103_ & new_n_n104_;
  assign new_n_n125_ = new_nd1_ & new_nn2_;
  assign new_n_n0_ = ~new_nm8_;
  assign new_nm3_ = new_n_n58_ & new_nt0_ & new_n_n75_;
  assign new_n_n367_ = new_nn2_ & new_n_n9_ & new_n_n8_ & new_ne1_;
  assign new_n_n341_ = new_n_n108_ & new_nj1_ & new_n_n58_;
  assign new_n_n324_ = new_n_n75_ & new_ni_ & new_n_n18_ & new_ng0_;
  assign new_nq4_ = new_n_n299_ | new_n_n298_ | new_n_n297_;
  assign new_n_n291_ = new_n_n75_ & new_n_n40_ & new_n_n30_ & new_n_n80_;
  assign new_nb5_ = new_n_n266_ | new_n_n265_ | new_n_n264_;
  assign new_ne5_ = new_n_n255_ | new_n_n254_ | new_n_n257_ | new_n_n256_ | new_n_n253_ | new_n_n252_ | new_n_n258_ | new_n_n251_;
  assign new_n_n219_ = new_n_n109_ & new_n_n55_ & new_n_n49_;
  assign new_n_n209_ = new_n_n52_ & new_nq2_ & new_n_n51_;
  assign new_n_n195_ = new_n_n111_ & new_nr2_ & new_n_n58_;
  assign new_n_n178_ = new_n_n75_ & new_nb1_ & new_nn1_;
  assign new_no5_ = new_n_n168_ | new_n_n169_;
  assign new_nc11_ = new_n_n145_ | new_n_n147_ | new_n_n146_ | new_n_n148_;
  assign new_ni11_ = new_n_n76_ | new_n_n77_ | new_ni0_;
  assign new_nc12_ = new_n_n108_ | new_n_n87_;
  assign new_nj13_ = new_n_n108_ | new_n_n98_;
  assign new_nw13_ = new_n_n132_ | new_nu2_;
  assign new_n_n126_ = new_nn2_ & new_ne1_;
  assign new_n_n1_ = ~new_nk8_;
  assign new_nn3_ = new_nb_ & new_n_n75_;
  assign new_n_n368_ = new_nv2_ & new_ng0_ & new_n_n7_;
  assign new_n_n332_ = new_n_n12_ & new_nk1_ & new_n_n58_;
  assign new_n_n331_ = new_nt0_ & new_n_n11_ & new_n_n58_;
  assign new_n_n299_ = new_n_n75_ & new_n_n41_ & new_nx1_;
  assign new_n_n292_ = new_ng0_ & new_n_n42_ & new_nu_ & new_n_n81_;
  assign new_n_n266_ = new_n_n75_ & new_n_n41_ & new_ni2_;
  assign new_n_n259_ = new_n_n43_ & new_n_n60_;
  assign new_n_n218_ = new_n_n111_ & new_n_n55_ & new_n_n49_;
  assign new_n_n210_ = new_n_n50_ & new_nq2_ & new_n_n51_;
  assign new_n_n185_ = new_nd1_ & new_n_n53_ & new_n_n58_ & new_n_n52_;
  assign new_n_n177_ = new_n_n75_ & new_ne1_ & new_nn1_ & new_n_n80_;
  assign new_n_n170_ = new_n_n59_ & new_n_n60_;
  assign new_n_n148_ = new_ne1_ & new_n_n80_;
  assign new_n_n141_ = new_n_n75_ & new_ne1_ & new_np1_ & new_n_n80_;
  assign new_nf12_ = new_n_n108_ | new_n_n88_;
  assign new_ng13_ = new_n_n108_ | new_n_n97_;
  assign new_n_n132_ = new_nb_ & new_n_n101_;
  assign new_na14_ = new_n_n124_ | new_n_n126_ | new_n_n125_ | new_nc1_;
  assign new_n_n2_ = ~new_nj8_;
  assign new_n_n370_ = new_nv2_ & new_ng0_ & new_n_n7_ & new_n_n58_;
  assign new_n_n361_ = new_no0_ & new_nf1_ & new_n_n58_;
  assign new_n_n352_ = new_nn2_ & new_nh1_ & new_n_n58_;
  assign new_nc4_ = new_n_n339_ | new_n_n359_ | new_n_n341_ | new_n_n340_ | new_n_n338_ | new_n_n337_ | new_n_n342_ | new_n_n336_;
  assign new_n_n333_ = new_nt0_ & new_nk1_ & new_n_n58_;
  assign new_ne4_ = new_n_n329_ | new_n_n330_;
  assign new_ni4_ = new_n_n323_ | new_n_n322_ | new_n_n321_;
  assign new_n_n315_ = new_n_n75_ & new_n_n40_ & new_n_n22_ & new_n_n80_;
  assign new_n_n307_ = new_ng0_ & new_n_n42_ & new_np_ & new_n_n81_;
  assign new_nv4_ = new_n_n284_ | new_n_n283_ | new_n_n282_;
  assign new_n_n276_ = new_n_n75_ & new_n_n40_ & new_n_n35_ & new_n_n80_;
  assign new_n_n268_ = new_ng0_ & new_n_n42_ & new_nc0_ & new_n_n81_;
  assign new_n_n260_ = new_n_n43_ & new_nk2_;
  assign new_n_n258_ = new_n_n104_ & new_nl2_ & new_n_n44_;
  assign new_n_n248_ = new_n_n102_ & new_nu2_ & new_n_n45_;
  assign new_nh5_ = new_n_n233_ | new_n_n232_ | new_n_n230_ | new_n_n229_ | new_n_n231_ | new_n_n237_ | new_n_n235_ | new_n_n234_ | new_n_n228_ | new_n_n236_ | new_n_n238_;
  assign new_n_n228_ = new_n_n55_ & new_n_n52_ & new_n_n48_;
  assign new_n_n213_ = new_n_n55_ & new_n_n52_ & new_n_n49_;
  assign new_n_n200_ = new_n_n111_ & new_n_n55_ & new_n_n51_;
  assign new_n_n190_ = new_n_n109_ & new_n_n53_ & new_n_n58_ & new_nd1_;
  assign new_n_n180_ = new_n_n75_ & new_nm0_ & new_nb1_;
  assign new_n_n171_ = new_n_n59_ & new_nk2_;
  assign new_n_n163_ = new_nm1_ & new_nh_;
  assign new_n_n156_ = new_n_n66_ & new_no2_;
  assign new_n_n150_ = new_n_n71_ & new_n_n73_ & new_nh0_ & new_n_n72_;
  assign new_nf11_ = new_n_n141_ | new_n_n143_ | new_n_n142_ | new_n_n144_;
  assign new_n_n137_ = new_n_n79_ & new_nv2_ & new_nm1_ & new_ng0_;
  assign new_n_n135_ = new_nv2_ & new_ng0_ & new_n_n81_ & new_nm1_;
  assign new_nr12_ = new_n_n108_ | new_n_n92_;
  assign new_n_n134_ = new_nu2_ & new_nk2_;
  assign new_nz13_ = new_n_n102_ | new_n_n103_ | new_nk2_;
  assign new_n_n113_ = new_nq2_ & new_n_n111_ & new_nr2_ & new_n_n112_;
  assign new_n_n102_ = ~new_nm2_;
  assign new_nx2_ = ~new_ng1_;
  assign new_nd3_ = new_n_n370_ | new_n_n3_;
  assign new_n_n360_ = new_n_n12_ & new_nf1_ & new_n_n58_;
  assign new_na4_ = new_n_n349_ | new_n_n359_ | new_n_n351_ | new_n_n350_ | new_n_n338_ | new_n_n348_ | new_n_n352_ | new_n_n336_;
  assign new_n_n342_ = new_nn2_ & new_nj1_ & new_n_n58_;
  assign new_n_n334_ = new_n_n108_ & new_nk1_ & new_n_n58_;
  assign new_n_n330_ = new_nl1_ & new_n_n58_;
  assign new_nh4_ = new_n_n135_ | new_n_n19_;
  assign new_nl4_ = new_n_n314_ | new_n_n313_ | new_n_n312_;
  assign new_n_n308_ = new_n_n75_ & new_n_n41_ & new_nu1_;
  assign new_n_n284_ = new_n_n75_ & new_n_n41_ & new_nc2_;
  assign new_n_n277_ = new_ng0_ & new_n_n42_ & new_nz_ & new_n_n81_;
  assign new_n_n267_ = new_n_n75_ & new_n_n40_ & new_n_n38_ & new_n_n80_;
  assign new_n_n261_ = new_n_n43_ & new_nu2_;
  assign new_n_n257_ = new_n_n104_ & new_nu2_ & new_n_n44_;
  assign new_n_n249_ = new_n_n103_ & new_nu2_ & new_n_n45_;
  assign new_n_n238_ = new_n_n109_ & new_no2_ & new_n_n48_;
  assign new_n_n229_ = new_nd1_ & new_n_n52_ & new_n_n48_;
  assign new_n_n204_ = new_n_n111_ & new_nd1_ & new_n_n51_;
  assign new_n_n199_ = new_n_n109_ & new_n_n55_ & new_n_n51_;
  assign new_n_n191_ = new_n_n111_ & new_n_n53_ & new_n_n58_ & new_ne1_;
  assign new_n_n179_ = new_n_n75_ & new_n_n108_ & new_nb1_;
  assign new_n_n172_ = new_n_n59_ & new_n_n103_;
  assign new_n_n168_ = new_n_n67_ & new_nv2_ & new_n_n62_;
  assign new_n_n155_ = new_n_n66_ & new_n_n109_;
  assign new_ng10_ = new_n_n150_ | new_ng0_ | new_nm1_ | new_n_n75_;
  assign new_n_n144_ = new_n_n75_ & new_nm0_ & new_n_n74_;
  assign new_n_n138_ = new_ni_ & new_nv2_ & new_nm1_ & new_ng0_;
  assign new_nn11_ = new_n_n108_ | new_n_n82_;
  assign new_no12_ = new_n_n108_ | new_n_n91_;
  assign new_n_n133_ = new_n_n101_ & new_nb_ & new_nk2_;
  assign new_n_n127_ = new_n_n102_ & new_n_n103_;
  assign new_n_n112_ = ~new_np2_;
  assign new_n_n103_ = ~new_nl2_;
  assign new_ny2_ = ~new_nh1_;
  assign new_n_n371_ = new_n_n75_ & new_n_n2_ & new_n_n1_ & new_ne1_;
  assign new_nq3_ = new_n_n75_ & new_nw0_;
  assign new_n_n359_ = new_nn2_ & new_n_n11_ & new_n_n58_;
  assign new_n_n350_ = new_nq0_ & new_nh1_ & new_n_n58_;
  assign new_n_n344_ = new_n_n12_ & new_ni1_ & new_n_n58_;
  assign new_n_n335_ = new_nn2_ & new_nk1_ & new_n_n58_;
  assign new_n_n329_ = new_n_n58_ & new_nn2_ & new_n_n13_ & new_ne1_;
  assign new_n_n322_ = new_ng0_ & new_nk_ & new_n_n42_ & new_n_n81_;
  assign new_n_n317_ = new_n_n75_ & new_n_n41_ & new_nr1_;
  assign new_nn4_ = new_n_n308_ | new_n_n307_ | new_n_n306_;
  assign new_nr4_ = new_n_n296_ | new_n_n295_ | new_n_n294_;
  assign new_n_n288_ = new_n_n75_ & new_n_n40_ & new_n_n31_ & new_n_n80_;
  assign new_n_n283_ = new_ng0_ & new_n_n42_ & new_nx_ & new_n_n81_;
  assign new_n_n275_ = new_n_n75_ & new_n_n41_ & new_nf2_;
  assign new_na5_ = new_n_n269_ | new_n_n268_ | new_n_n267_;
  assign new_nd5_ = new_n_n261_ | new_n_n260_ | new_n_n259_;
  assign new_n_n256_ = new_n_n103_ & new_nu2_ & new_n_n44_;
  assign new_n_n246_ = new_n_n102_ & new_n_n60_ & new_n_n45_;
  assign new_n_n240_ = new_n_n47_ & new_nd1_;
  assign new_n_n230_ = new_ne1_ & new_n_n52_ & new_n_n48_;
  assign new_n_n215_ = new_ne1_ & new_n_n52_ & new_n_n49_;
  assign new_n_n205_ = new_n_n52_ & new_ne1_ & new_n_n51_;
  assign new_n_n198_ = new_n_n50_ & new_n_n55_ & new_n_n51_;
  assign new_n_n188_ = new_n_n109_ & new_n_n53_ & new_n_n58_ & new_n_n55_;
  assign new_n_n181_ = new_n_n55_ & new_n_n53_ & new_n_n58_ & new_n_n54_;
  assign new_n_n173_ = new_n_n59_ & new_n_n102_;
  assign new_nj8_ = new_n_n109_ | new_np2_ | new_no2_ | new_n_n68_;
  assign new_n_n161_ = new_nm1_ & new_n_n79_;
  assign new_n_n151_ = new_n_n76_ & new_n_n75_;
  assign new_n_n145_ = new_nv2_ & new_nh_ & new_nm1_ & new_ng0_;
  assign new_n_n139_ = new_nh_ & new_nv2_ & new_nm1_ & new_ng0_;
  assign new_nq11_ = new_n_n108_ | new_n_n83_;
  assign new_nx12_ = new_n_n108_ | new_n_n94_;
  assign new_nu13_ = new_n_n106_ | new_nu0_;
  assign new_n_n128_ = new_n_n102_ & new_n_n104_;
  assign new_nb14_ = new_ne1_ | new_nd1_ | new_n_n123_;
  assign new_n_n117_ = new_n_n105_ & new_n_n112_;
  assign new_nz2_ = ~new_ni1_;
  assign new_n_n372_ = new_n_n75_ & new_ns2_ & new_n_n0_;
  assign new_n_n366_ = new_ne1_ & new_n_n58_;
  assign new_n_n358_ = new_no0_ & new_n_n11_ & new_n_n58_;
  assign new_n_n351_ = new_n_n108_ & new_nh1_ & new_n_n58_;
  assign new_n_n343_ = new_nr0_ & new_n_n11_ & new_n_n58_;
  assign new_nd4_ = new_n_n332_ | new_n_n359_ | new_n_n334_ | new_n_n333_ | new_n_n338_ | new_n_n331_ | new_n_n335_ | new_n_n336_;
  assign new_nf4_ = new_n_n327_ | new_n_n328_;
  assign new_n_n323_ = new_n_n75_ & new_np1_ & new_n_n41_;
  assign new_n_n316_ = new_ng0_ & new_n_n42_ & new_nm_ & new_n_n81_;
  assign new_n_n309_ = new_n_n75_ & new_n_n40_ & new_n_n24_ & new_n_n80_;
  assign new_n_n296_ = new_n_n75_ & new_n_n41_ & new_ny1_;
  assign new_n_n289_ = new_ng0_ & new_n_n42_ & new_nv_ & new_n_n81_;
  assign new_n_n282_ = new_n_n75_ & new_n_n40_ & new_n_n33_ & new_n_n80_;
  assign new_ny4_ = new_n_n275_ | new_n_n274_ | new_n_n273_;
  assign new_n_n269_ = new_n_n75_ & new_n_n41_ & new_nh2_;
  assign new_n_n262_ = new_ng0_ & new_n_n42_ & new_n_n81_ & new_ne0_;
  assign new_n_n255_ = new_n_n104_ & new_n_n60_ & new_n_n44_;
  assign new_n_n247_ = new_n_n103_ & new_n_n60_ & new_n_n45_;
  assign new_n_n239_ = new_n_n47_ & new_n_n55_;
  assign new_n_n231_ = new_no2_ & new_n_n52_ & new_n_n48_;
  assign new_n_n214_ = new_nd1_ & new_n_n52_ & new_n_n49_;
  assign new_n_n206_ = new_n_n50_ & new_ne1_ & new_n_n51_;
  assign new_n_n197_ = new_n_n52_ & new_n_n55_ & new_n_n51_;
  assign new_n_n189_ = new_n_n111_ & new_n_n53_ & new_n_n58_ & new_nd1_;
  assign new_nl5_ = new_n_n177_ | new_n_n179_ | new_n_n178_ | new_n_n180_;
  assign new_nn5_ = new_n_n170_ | new_n_n172_ | new_n_n171_ | new_n_n173_;
  assign new_nk8_ = new_n_n165_ | new_n_n167_ | new_n_n166_;
  assign new_n_n162_ = new_nm1_ & new_ni_;
  assign new_nk9_ = new_n_n153_ | new_n_n155_ | new_n_n154_ | new_n_n156_;
  assign new_ne11_ = new_nh0_ & new_n_n72_ & new_n_n71_ & new_n_n73_;
  assign new_n_n140_ = new_ng_ & new_nv2_ & new_nm1_ & new_ng0_;
  assign new_nt11_ = new_n_n108_ | new_n_n84_;
  assign new_nu12_ = new_n_n108_ | new_n_n93_;
  assign new_nv13_ = new_nc1_ | new_n_n134_ | new_n_n133_;
  assign new_n_n129_ = new_nl2_ & new_n_n104_;
  assign new_n_n123_ = new_n_n104_ & new_nl2_ & new_nm2_;
  assign new_n_n118_ = new_n_n105_ & new_n_n111_;
  assign new_na3_ = ~new_nj1_;
  assign new_n_n88_ = ~new_nx1_;
  assign new_n_n77_ = ~new_nm1_;
  assign new_n_n66_ = ~new_nn0_;
  assign new_n_n55_ = ~new_nz13_;
  assign new_n_n44_ = ~new_nx13_;
  assign new_n_n89_ = ~new_ny1_;
  assign new_n_n76_ = ~new_nv2_;
  assign new_n_n67_ = ~new_nf0_;
  assign new_n_n54_ = ~new_ng14_;
  assign new_n_n45_ = ~new_ny13_;
  assign new_n_n90_ = ~new_nz1_;
  assign new_n_n75_ = ~new_ni0_;
  assign new_n_n64_ = ~new_no8_;
  assign new_n_n57_ = ~new_ns2_;
  assign new_n_n46_ = ~new_nw13_;
  assign new_n_n91_ = ~new_na2_;
  assign new_n_n74_ = ~new_no1_;
  assign new_n_n65_ = ~new_nk0_;
  assign new_n_n56_ = ~new_nl1_;
  assign new_n_n47_ = ~new_na14_;
  assign new_nw2_ = ~new_nf1_;
  assign new_n_n92_ = ~new_nb2_;
  assign new_n_n37_ = ~new_nj13_;
  assign new_n_n26_ = ~new_nc12_;
  assign new_n_n15_ = ~new_nc11_;
  assign new_n_n4_ = ~new_ni9_;
  assign new_n_n93_ = ~new_nc2_;
  assign new_n_n36_ = ~new_ng13_;
  assign new_n_n27_ = ~new_nf12_;
  assign new_n_n14_ = ~new_nu10_;
  assign new_n_n5_ = ~new_nk9_;
  assign new_n_n35_ = ~new_nd13_;
  assign new_n_n24_ = ~new_nw11_;
  assign new_n_n17_ = ~new_ny10_;
  assign new_n_n6_ = ~new_nf10_;
  assign new_n_n34_ = ~new_na13_;
  assign new_n_n25_ = ~new_nz11_;
  assign new_n_n16_ = ~new_nz10_;
  assign new_n_n7_ = ~new_nw8_;
  assign new_n_n63_ = ~new_nt2_;
  assign new_n_n52_ = ~new_nb14_;
  assign new_n_n41_ = ~new_nl11_;
  assign new_n_n30_ = ~new_no12_;
  assign new_n_n19_ = ~new_nf11_;
  assign new_n_n8_ = ~new_ne10_;
  assign new_n_n62_ = ~new_nv10_;
  assign new_n_n53_ = ~new_nh14_;
  assign new_n_n40_ = ~new_nk11_;
  assign new_n_n31_ = ~new_nr12_;
  assign new_n_n18_ = ~new_na11_;
  assign new_n_n9_ = ~new_nd10_;
  assign new_n_n83_ = ~new_ns1_;
  assign new_n_n72_ = ~new_nh_;
  assign new_n_n39_ = ~new_np13_;
  assign new_n_n28_ = ~new_ni12_;
  assign new_n_n21_ = ~new_nn11_;
  assign new_n_n10_ = ~new_ng10_;
  assign new_n_n82_ = ~new_nr1_;
  assign new_n_n73_ = ~new_ni_;
  assign new_n_n38_ = ~new_nm13_;
  assign new_n_n29_ = ~new_nl12_;
  assign new_n_n20_ = ~new_nj11_;
  assign new_n_n11_ = ~new_nn10_;
  assign new_n_n84_ = ~new_nt1_;
  assign new_n_n81_ = ~new_ne11_;
  assign new_n_n70_ = ~new_nx10_;
  assign new_n_n59_ = ~new_nj14_;
  assign new_n_n48_ = ~new_nc14_;
  assign new_n_n23_ = ~new_nt11_;
  assign new_n_n12_ = ~new_nl10_;
  assign new_n_n85_ = ~new_nu1_;
  assign new_n_n80_ = ~new_nm0_;
  assign new_n_n71_ = ~new_ng_;
  assign new_n_n58_ = ~new_nc1_;
  assign new_n_n49_ = ~new_nd14_;
  assign new_n_n22_ = ~new_nq11_;
  assign new_n_n13_ = ~new_nf9_;
  assign new_n_n86_ = ~new_nv1_;
  assign new_n_n79_ = ~new_nh0_;
  assign new_n_n68_ = ~new_nr2_;
  assign new_n_n61_ = ~new_nk14_;
  assign new_n_n50_ = ~new_ne14_;
  assign new_n_n43_ = ~new_nv13_;
  assign new_n_n32_ = ~new_nu12_;
  assign new_n_n87_ = ~new_nw1_;
  assign new_n_n78_ = ~new_nq1_;
  assign new_n_n69_ = ~new_nl9_;
  assign new_n_n60_ = ~new_nu13_;
  assign new_n_n51_ = ~new_nf14_;
  assign new_n_n42_ = ~new_ni11_;
  assign new_n_n33_ = ~new_nx12_;
endmodule


