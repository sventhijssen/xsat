// Benchmark "top" written by ABC on Fri Mar 31 12:13:06 2023

module top ( 
    pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1, pf4, pr,
    pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0, pf3,
    pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, pk3, pl4, px, ph1, pi0, pj3, pk2, pm4, py, ph2, pi3, pj0,
    pk1, pn4, pz, ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pi4, pl1,
    pm0, pn3, po2, pj4, pl2, pm3, pn0, po1, pk4, pl3, pm2, pn1, po0, pp0,
    pq1, pr2, ps3, pa, pp1, pq0, pr3, ps2, pb, pp2, pq3, ps1, pc, pp3, pq2,
    pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1, pu0, pv3, pw2, pf, pt2, pu3,
    pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1, py0, pz3,
    pj, px2, py3, pz0, pk, px3, py2, pz1, pl, pm, pn, po,
    pe5, pf6, pg7, ph8, pi9, pd5, pf7, pg6, ph9, pi8, pd6, pe7, pg5, pj8,
    pk9, pd7, pe6, pf5, pj9, pk8, pa5, pb6, pc7, pl8, pm9, pb7, pc6, pl9,
    pm8, pa7, pc5, pn8, po9, pa6, pb5, pn9, po8, pa9, pm5, pn6, po7, pa8,
    pl5, pn7, po6, pb8, pc9, pl6, pm7, po5, pb9, pc8, pl7, pm6, pn5, po4,
    pd8, pe9, pi5, pj6, pk7, pd9, pe8, ph5, pj7, pk6, pf8, pg9, ph6, pi7,
    pk5, pf9, pg8, ph7, pi6, pj5, pt4, pu5, pv6, pw7, px8, pt5, pu4, pv7,
    pw6, py8, pt6, pu7, pv4, pw5, pz8, pt7, pu6, pv5, pw4, pp4, pq5, pr6,
    ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7, pq6, pr5, ps4, pp8,
    pq9, pp9, pq8, pr8, ps9, pr9, ps8, pt8, pu9, px4, py5, pz6, pt9, pu8,
    px5, py4, pz7, pv8, pw9, px6, py7, pz4, pv9, pw8, px7, py6, pz5  );
  input  pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1,
    pf4, pr, pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0,
    pf3, pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw,
    ph0, pi1, pj2, pk3, pl4, px, ph1, pi0, pj3, pk2, pm4, py, ph2, pi3,
    pj0, pk1, pn4, pz, ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pi4,
    pl1, pm0, pn3, po2, pj4, pl2, pm3, pn0, po1, pk4, pl3, pm2, pn1, po0,
    pp0, pq1, pr2, ps3, pa, pp1, pq0, pr3, ps2, pb, pp2, pq3, ps1, pc, pp3,
    pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1, pu0, pv3, pw2, pf, pt2,
    pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1, py0,
    pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, pm, pn, po;
  output pe5, pf6, pg7, ph8, pi9, pd5, pf7, pg6, ph9, pi8, pd6, pe7, pg5, pj8,
    pk9, pd7, pe6, pf5, pj9, pk8, pa5, pb6, pc7, pl8, pm9, pb7, pc6, pl9,
    pm8, pa7, pc5, pn8, po9, pa6, pb5, pn9, po8, pa9, pm5, pn6, po7, pa8,
    pl5, pn7, po6, pb8, pc9, pl6, pm7, po5, pb9, pc8, pl7, pm6, pn5, po4,
    pd8, pe9, pi5, pj6, pk7, pd9, pe8, ph5, pj7, pk6, pf8, pg9, ph6, pi7,
    pk5, pf9, pg8, ph7, pi6, pj5, pt4, pu5, pv6, pw7, px8, pt5, pu4, pv7,
    pw6, py8, pt6, pu7, pv4, pw5, pz8, pt7, pu6, pv5, pw4, pp4, pq5, pr6,
    ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7, pq6, pr5, ps4, pp8,
    pq9, pp9, pq8, pr8, ps9, pr9, ps8, pt8, pu9, px4, py5, pz6, pt9, pu8,
    px5, py4, pz7, pv8, pw9, px6, py7, pz4, pv9, pw8, px7, py6, pz5;
  wire new_na1_, new_nb2_, new_nc3_, new_nd4_, new_np_, new_na0_, new_nb3_,
    new_nc2_, new_ne4_, new_nq_, new_na3_, new_nb0_, new_nc1_, new_nf4_,
    new_nr_, new_na2_, new_nb1_, new_nc0_, new_ng4_, new_ns_, new_nd0_,
    new_ne1_, new_nf2_, new_ng3_, new_nt_, new_na4_, new_nd1_, new_ne0_,
    new_nf3_, new_ng2_, new_nu_, new_nb4_, new_nd2_, new_ne3_, new_nf0_,
    new_ng1_, new_nv_, new_nc4_, new_nd3_, new_ne2_, new_nf1_, new_ng0_,
    new_nw_, new_nh0_, new_ni1_, new_nj2_, new_nk3_, new_nl4_, new_nx_,
    new_nh1_, new_ni0_, new_nj3_, new_nk2_, new_nm4_, new_ny_, new_nh2_,
    new_ni3_, new_nj0_, new_nk1_, new_nn4_, new_nz_, new_nh3_, new_ni2_,
    new_nj1_, new_nk0_, new_nh4_, new_nl0_, new_nm1_, new_nn2_, new_no3_,
    new_ni4_, new_nl1_, new_nm0_, new_nn3_, new_no2_, new_nj4_, new_nl2_,
    new_nm3_, new_nn0_, new_no1_, new_nk4_, new_nl3_, new_nm2_, new_nn1_,
    new_no0_, new_np0_, new_nq1_, new_nr2_, new_ns3_, new_na_, new_np1_,
    new_nq0_, new_nr3_, new_ns2_, new_nb_, new_np2_, new_nq3_, new_ns1_,
    new_nc_, new_np3_, new_nq2_, new_nr1_, new_ns0_, new_nd_, new_nt0_,
    new_nu1_, new_nv2_, new_nw3_, new_ne_, new_nt1_, new_nu0_, new_nv3_,
    new_nw2_, new_nf_, new_nt2_, new_nu3_, new_nv0_, new_nw1_, new_ng_,
    new_nt3_, new_nu2_, new_nv1_, new_nw0_, new_nh_, new_nx0_, new_ny1_,
    new_nz2_, new_ni_, new_nx1_, new_ny0_, new_nz3_, new_nj_, new_nx2_,
    new_ny3_, new_nz0_, new_nk_, new_nx3_, new_ny2_, new_nz1_, new_nl_,
    new_nm_, new_nn_, new_no_, new_n_n1007_, new_n_n997_, new_n_n920_,
    new_n_n910_, new_n_n900_, new_n_n890_, new_n_n880_, new_n_n833_,
    new_nw7_, new_nh8_, new_n_n819_, new_np8_, new_n_n804_, new_n_n797_,
    new_na9_, new_n_n770_, new_nq9_, new_nv9_, new_no15_, new_n_n749_,
    new_nm16_, new_na17_, new_nl17_, new_nx17_, new_nm19_, new_n_n712_,
    new_ni20_, new_nu20_, new_n_n699_, new_nj21_, new_n_n687_, new_na22_,
    new_n_n676_, new_nt22_, new_n_n663_, new_ni23_, new_n_n630_, new_nl24_,
    new_n_n616_, new_nw24_, new_nd25_, new_n_n600_, new_nr25_, new_ng27_,
    new_nw27_, new_n_n590_, new_nm28_, new_nu28_, new_nx28_, new_nj29_,
    new_n_n559_, new_na30_, new_nl30_, new_n_n544_, new_ni31_, new_n_n541_,
    new_na32_, new_nl32_, new_n_n530_, new_nx32_, new_nh33_, new_nl33_,
    new_n_n507_, new_n_n501_, new_nx33_, new_n_n486_, new_nk34_, new_nw34_,
    new_n_n475_, new_n_n469_, new_nl35_, new_n_n457_, new_nj6_,
    new_n_n439_, new_n_n428_, new_n_n417_, new_n_n406_, new_n_n396_,
    new_no4_, new_n_n364_, new_n_n353_, new_n_n342_, new_n_n331_,
    new_n_n320_, new_n_n309_, new_n_n298_, new_n_n287_, new_n_n254_,
    new_n_n243_, new_n_n232_, new_n_n221_, new_n_n210_, new_n_n199_,
    new_n_n188_, new_n_n144_, new_n_n133_, new_n_n122_, new_n_n111_,
    new_n_n100_, new_n_n89_, new_n_n1006_, new_n_n998_, new_n_n919_,
    new_n_n911_, new_n_n899_, new_n_n891_, new_n_n871_, new_n_n832_,
    new_nv7_, new_ni8_, new_nl8_, new_n_n811_, new_n_n805_, new_n_n796_,
    new_n_n790_, new_nh9_, new_n_n763_, new_nu9_, new_n_n753_, new_n_n750_,
    new_np16_, new_n_n742_, new_nn17_, new_nv17_, new_n_n716_, new_nw19_,
    new_nk20_, new_ns20_, new_nf21_, new_n_n692_, new_ns21_, new_nz21_,
    new_n_n675_, new_n_n670_, new_n_n662_, new_n_n657_, new_n_n629_,
    new_n_n623_, new_n_n615_, new_n_n609_, new_ne25_, new_n_n601_,
    new_nx25_, new_nh27_, new_nv27_, new_n_n589_, new_n_n582_, new_n_n576_,
    new_nw28_, new_n_n565_, new_n_n560_, new_nb30_, new_nk30_, new_nv30_,
    new_nh31_, new_nr31_, new_nz31_, new_nm32_, new_n_n531_, new_n_n522_,
    new_n_n521_, new_n_n515_, new_np33_, new_nt33_, new_n_n493_,
    new_n_n487_, new_nl34_, new_nv34_, new_n_n474_, new_nh35_, new_n_n468_,
    new_n_n456_, new_n_n447_, new_n_n438_, new_n_n429_, new_n_n416_,
    new_n_n407_, new_n_n395_, new_n_n386_, new_n_n363_, new_n_n354_,
    new_n_n341_, new_n_n332_, new_n_n319_, new_n_n310_, new_n_n297_,
    new_n_n288_, new_n_n264_, new_n_n242_, new_n_n233_, new_n_n220_,
    new_n_n211_, new_n_n198_, new_n_n189_, new_n_n143_, new_n_n134_,
    new_n_n121_, new_n_n112_, new_n_n99_, new_n_n90_, new_ny4_,
    new_n_n1009_, new_n_n999_, new_n_n922_, new_n_n912_, new_n_n898_,
    new_n_n882_, new_n_n872_, new_ns7_, new_nu7_, new_n_n825_, new_nm8_,
    new_n_n813_, new_ns8_, new_nd9_, new_n_n776_, new_n_n762_, new_n_n756_,
    new_nl15_, new_nb16_, new_n_n745_, new_nd17_, new_nj17_, new_n_n734_,
    new_ns18_, new_n_n720_, new_n_n707_, new_nv20_, new_nc21_, new_n_n693_,
    new_n_n689_, new_n_n682_, new_nm22_, new_n_n668_, new_na23_,
    new_n_n658_, new_n_n632_, new_n_n624_, new_ns24_, new_ny24_,
    new_n_n607_, new_ni25_, new_nm26_, new_nd27_, new_nt27_, new_n_n588_,
    new_n_n581_, new_n_n578_, new_nv28_, new_n_n554_, new_nx29_, new_nj30_,
    new_nw30_, new_n_n542_, new_nq31_, new_ny31_, new_nn32_, new_nw32_,
    new_ne33_, new_nq33_, new_nu33_, new_n_n495_, new_na34_, new_nm34_,
    new_n_n483_, new_n_n476_, new_ng35_, new_n_n455_, new_n_n446_,
    new_n_n441_, new_n_n430_, new_n_n415_, new_n_n404_, new_n_n398_,
    new_n_n387_, new_n_n362_, new_n_n351_, new_n_n344_, new_n_n333_,
    new_n_n318_, new_n_n307_, new_n_n300_, new_n_n289_, new_n_n263_,
    new_n_n252_, new_n_n234_, new_n_n219_, new_n_n208_, new_n_n201_,
    new_n_n190_, new_n_n164_, new_n_n153_, new_n_n120_, new_n_n109_,
    new_n_n102_, new_n_n91_, new_n_n1072_, new_n_n1008_, new_n_n1000_,
    new_n_n921_, new_n_n913_, new_n_n889_, new_n_n881_, new_n_n873_,
    new_n_n834_, new_nt7_, new_n_n824_, new_n_n818_, new_n_n812_,
    new_n_n806_, new_n_n783_, new_n_n777_, new_nr9_, new_n_n757_,
    new_nm15_, new_nz15_, new_nr16_, new_nb17_, new_n_n738_, new_nt17_,
    new_n_n724_, new_nc19_, new_nl20_, new_n_n703_, new_ne21_, new_n_n694_,
    new_n_n688_, new_n_n683_, new_n_n674_, new_n_n669_, new_n_n664_,
    new_n_n659_, new_n_n631_, new_n_n625_, new_n_n614_, new_nx24_,
    new_n_n606_, new_nh25_, new_nb27_, new_ne27_, new_ns27_, new_n_n587_,
    new_nn28_, new_n_n577_, new_n_n569_, new_n_n553_, new_nw29_, new_ny29_,
    new_nx30_, new_nj31_, new_nz29_, new_nw31_, new_n_n529_, new_n_n526_,
    new_n_n523_, new_n_n506_, new_n_n500_, new_n_n494_, new_n_n488_,
    new_nn34_, new_nx34_, new_nb35_, new_nf35_, new_n_n454_, new_nk6_,
    new_n_n440_, new_n_n431_, new_n_n414_, new_n_n405_, new_n_n397_,
    new_n_n388_, new_n_n361_, new_n_n352_, new_n_n343_, new_n_n334_,
    new_n_n317_, new_n_n308_, new_n_n299_, new_n_n290_, new_n_n262_,
    new_n_n253_, new_n_n244_, new_n_n218_, new_n_n209_, new_n_n200_,
    new_n_n191_, new_n_n163_, new_n_n154_, new_n_n119_, new_n_n110_,
    new_n_n101_, new_n_n92_, new_n_n1081_, new_n_n1073_, new_n_n1011_,
    new_n_n1001_, new_n_n924_, new_n_n914_, new_n_n864_, new_n_n854_,
    new_n_n844_, new_nj8_, new_n_n816_, new_nv8_, new_n_n792_, new_n_n785_,
    new_ng9_, new_n_n761_, new_ng15_, new_nw15_, new_n_n748_, new_nh16_,
    new_n_n744_, new_ni17_, new_n_n735_, new_nu18_, new_ng19_, new_n_n715_,
    new_nb20_, new_na21_, new_ni21_, new_n_n686_, new_nf22_, new_n_n677_,
    new_no22_, new_n_n666_, new_nh23_, new_n_n628_, new_no24_, new_n_n618_,
    new_nt24_, new_nb25_, new_ng25_, new_nm27_, new_nc28_, new_nh28_,
    new_n_n585_, new_nr28_, new_n_n570_, new_nd30_, new_no30_, new_n_n543_,
    new_no31_, new_nv31_, new_n_n519_, new_nm33_, new_n_n496_, new_n_n489_,
    new_n_n465_, new_np35_, new_n_n432_, new_n_n413_, new_n_n382_,
    new_n_n371_, new_n_n316_, new_n_n305_, new_n_n283_, new_n_n272_,
    new_n_n217_, new_n_n206_, new_n_n195_, new_n_n184_, new_n_n173_,
    new_n_n118_, new_n_n107_, new_n_n96_, new_n_n85_, new_n_n9_,
    new_n_n1080_, new_na5_, new_n_n1010_, new_n_n1002_, new_n_n923_,
    new_n_n915_, new_n_n863_, new_n_n855_, new_n_n835_, new_n_n823_,
    new_n_n817_, new_n_n799_, new_n_n793_, new_n_n784_, new_n_n778_,
    new_n_n760_, new_nw9_, new_n_n751_, new_nf16_, new_nj16_, new_nv16_,
    new_n_n739_, new_ns17_, new_nw18_, new_ne19_, new_nr19_, new_n_n711_,
    new_n_n700_, new_n_n695_, new_n_n685_, new_n_n680_, new_ng22_,
    new_nn22_, new_n_n665_, new_n_n660_, new_n_n627_, new_n_n621_,
    new_n_n617_, new_n_n611_, new_nc25_, new_nf25_, new_nn27_, new_nb28_,
    new_ni28_, new_nl28_, new_ns28_, new_n_n571_, new_ne30_, new_nn30_,
    new_nt30_, new_np31_, new_nu31_, new_n_n518_, new_n_n512_, new_nw33_,
    new_nz33_, new_ni35_, new_no35_, new_nl6_, new_n_n403_, new_n_n381_,
    new_n_n372_, new_n_n315_, new_n_n306_, new_n_n282_, new_n_n273_,
    new_n_n216_, new_n_n207_, new_n_n185_, new_n_n183_, new_n_n174_,
    new_n_n117_, new_n_n108_, new_n_n95_, new_n_n86_, new_nx4_,
    new_n_n1074_, new_n_n1013_, new_n_n1003_, new_nj7_, new_n_n862_,
    new_n_n846_, new_n_n836_, new_n_n810_, new_n_n803_, new_n_n798_,
    new_n_n791_, new_n_n786_, new_n_n779_, new_ns9_, new_n_n754_,
    new_n_n752_, new_nd16_, new_nl16_, new_n_n743_, new_n_n740_, new_nq17_,
    new_n_n723_, new_nh19_, new_no19_, new_na20_, new_ng20_, new_n_n704_,
    new_nt21_, new_n_n681_, new_nh22_, new_n_n671_, new_nv22_, new_n_n661_,
    new_nh24_, new_n_n622_, new_np24_, new_n_n610_, new_n_n608_,
    new_n_n602_, new_nj27_, new_nz27_, new_nj28_, new_n_n583_, new_n_n579_,
    new_n_n572_, new_n_n547_, new_nm30_, new_nu30_, new_nf31_, new_n_n539_,
    new_n_n520_, new_n_n513_, new_n_n509_, new_ns33_, new_n_n467_,
    new_nn35_, new_n_n448_, new_n_n394_, new_n_n384_, new_n_n373_,
    new_n_n296_, new_n_n285_, new_n_n274_, new_n_n215_, new_n_n197_,
    new_n_n186_, new_n_n116_, new_n_n105_, new_n_n98_, new_n_n87_,
    new_n_n1082_, new_n_n1075_, new_n_n1012_, new_n_n1004_, new_ni7_,
    new_n_n853_, new_n_n845_, new_n_n837_, new_nq8_, new_nt8_, new_nw8_,
    new_nz8_, new_nc9_, new_nf9_, new_n_n759_, new_n_n755_, new_nt15_,
    new_nc16_, new_n_n746_, new_nx16_, new_ng17_, new_n_n736_, new_nx18_,
    new_n_n719_, new_nq19_, new_ny19_, new_n_n708_, new_nq20_, new_nx21_,
    new_ne22_, new_nl22_, new_ns22_, new_nz22_, new_ng23_, new_ni24_,
    new_nm24_, new_nq24_, new_nu24_, new_na25_, new_n_n603_, new_nk27_,
    new_ny27_, new_n_n591_, new_n_n584_, new_nq28_, new_n_n573_, new_nc30_,
    new_n_n546_, new_n_n545_, new_ne31_, new_nn31_, new_ni33_, new_n_n514_,
    new_n_n508_, new_n_n502_, new_n_n466_, new_nm35_, new_n_n458_,
    new_n_n385_, new_n_n383_, new_n_n374_, new_n_n295_, new_n_n286_,
    new_n_n284_, new_n_n205_, new_n_n196_, new_n_n187_, new_n_n115_,
    new_n_n106_, new_n_n97_, new_n_n88_, new_nc5_, new_nk5_, new_n_n1057_,
    new_n_n1050_, new_n_n1041_, new_n_n995_, new_n_n985_, new_n_n975_,
    new_n_n965_, new_n_n955_, new_n_n945_, new_n_n935_, new_n_n925_,
    new_nl7_, new_n_n888_, new_n_n878_, new_n_n868_, new_n_n858_,
    new_n_n848_, new_n_n838_, new_n_n802_, new_n_n795_, new_nb9_,
    new_n_n780_, new_n_n772_, new_np9_, new_no17_, new_n_n731_, new_nn18_,
    new_n_n655_, new_nr23_, new_n_n643_, new_n_n635_, new_n_n599_,
    new_n_n595_, new_nd26_, new_nu26_, new_nb29_, new_nk29_, new_n_n556_,
    new_nt29_, new_nh30_, new_n_n536_, new_nr32_, new_ny32_, new_nk33_,
    new_no33_, new_n_n482_, new_n_n472_, new_n_n463_, new_n_n460_,
    new_n_n449_, new_n_n393_, new_n_n378_, new_n_n367_, new_n_n356_,
    new_n_n345_, new_n_n279_, new_n_n268_, new_n_n257_, new_n_n246_,
    new_n_n235_, new_n_n180_, new_n_n169_, new_n_n158_, new_n_n147_,
    new_n_n136_, new_n_n125_, new_n_n5_, new_n_n1067_, new_nj5_, new_no6_,
    new_n_n1051_, new_n_n1033_, new_n_n994_, new_n_n986_, new_n_n974_,
    new_n_n966_, new_n_n954_, new_n_n946_, new_n_n934_, new_n_n926_,
    new_nk7_, new_n_n887_, new_n_n879_, new_n_n867_, new_n_n859_,
    new_n_n847_, new_n_n839_, new_nu8_, new_nx8_, new_n_n787_, new_n_n781_,
    new_nl9_, new_n_n766_, new_ne17_, new_nd18_, new_n_n727_, new_nn23_,
    new_n_n649_, new_n_n642_, new_n_n636_, new_nl25_, new_n_n596_,
    new_nf26_, new_ns26_, new_nd29_, new_n_n564_, new_n_n555_, new_n_n550_,
    new_nr30_, new_nd32_, new_n_n528_, new_n_n524_, new_n_n516_,
    new_n_n510_, new_n_n481_, new_n_n473_, new_n_n462_, new_n_n461_,
    new_ni6_, new_n_n402_, new_n_n377_, new_n_n368_, new_n_n355_,
    new_n_n346_, new_n_n278_, new_n_n269_, new_n_n256_, new_n_n247_,
    new_n_n225_, new_n_n179_, new_n_n170_, new_n_n157_, new_n_n148_,
    new_n_n135_, new_n_n126_, new_n_n6_, new_n_n1066_, new_nw5_, new_nn6_,
    new_n_n1052_, new_n_n1024_, new_n_n993_, new_n_n983_, new_n_n977_,
    new_n_n967_, new_n_n953_, new_n_n943_, new_n_n937_, new_n_n927_,
    new_n_n906_, new_n_n896_, new_nn7_, new_n_n866_, new_n_n856_,
    new_n_n850_, new_n_n840_, new_n_n827_, new_nc8_, new_n_n801_, new_ny8_,
    new_n_n789_, new_ne9_, new_nk9_, new_no9_, new_nu16_, new_na18_,
    new_nm18_, new_n_n654_, new_nt23_, new_ny23_, new_n_n637_, new_nk24_,
    new_n_n598_, new_n_n594_, new_na26_, new_nr26_, new_np27_, new_nf28_,
    new_ne29_, new_nm29_, new_n_n558_, new_n_n551_, new_nf30_, new_nq30_,
    new_ne32_, new_n_n534_, new_n_n525_, new_n_n517_, new_n_n511_,
    new_nf34_, new_np34_, new_nj35_, new_nr35_, new_n_n433_, new_n_n412_,
    new_n_n380_, new_n_n369_, new_n_n336_, new_n_n325_, new_n_n281_,
    new_n_n270_, new_n_n255_, new_n_n237_, new_n_n226_, new_n_n182_,
    new_n_n171_, new_n_n156_, new_n_n145_, new_n_n138_, new_n_n127_,
    new_n_n7_, new_n_n1065_, new_nl5_, new_n_n1058_, new_n_n1053_,
    new_n_n1015_, new_n_n992_, new_n_n984_, new_n_n976_, new_n_n968_,
    new_n_n952_, new_n_n944_, new_n_n936_, new_n_n928_, new_n_n905_,
    new_n_n897_, new_nm7_, new_n_n865_, new_n_n857_, new_n_n849_,
    new_n_n841_, new_n_n826_, new_nb8_, new_n_n800_, new_n_n794_,
    new_n_n788_, new_n_n782_, new_n_n773_, new_n_n767_, new_ng16_,
    new_nc18_, new_nk18_, new_n_n653_, new_ns23_, new_n_n644_, new_n_n638_,
    new_n_n620_, new_nm25_, new_ns25_, new_nc26_, new_np26_, new_nq27_,
    new_ne28_, new_n_n567_, new_nl29_, new_n_n557_, new_n_n552_, new_ng30_,
    new_np30_, new_nf32_, new_n_n535_, new_nq32_, new_nj33_, new_nn33_,
    new_ng34_, new_no34_, new_n_n464_, new_nq35_, new_n_n423_, new_n_n422_,
    new_n_n379_, new_n_n370_, new_n_n335_, new_n_n326_, new_n_n280_,
    new_n_n271_, new_n_n245_, new_n_n236_, new_n_n227_, new_n_n181_,
    new_n_n172_, new_n_n155_, new_n_n146_, new_n_n137_, new_n_n128_,
    new_n_n8_, new_n_n1103_, new_nd5_, new_n_n1044_, new_n_n1035_,
    new_n_n1026_, new_n_n1016_, new_n_n991_, new_n_n981_, new_n_n971_,
    new_n_n961_, new_n_n959_, new_n_n949_, new_n_n939_, new_n_n929_,
    new_n_n916_, new_n_n904_, new_n_n894_, new_n_n884_, new_n_n874_,
    new_np7_, new_n_n852_, new_n_n842_, new_n_n829_, new_na8_, new_nd8_,
    new_nk8_, new_n_n814_, new_n_n807_, new_n_n774_, new_nn9_, new_ny15_,
    new_ny17_, new_n_n728_, new_n_n652_, new_n_n648_, new_na24_,
    new_n_n633_, new_n_n613_, new_nn25_, new_n_n592_, new_nj26_, new_na27_,
    new_n_n586_, new_np28_, new_n_n566_, new_n_n563_, new_nq29_, new_nv29_,
    new_nb31_, new_nl31_, new_n_n540_, new_ni32_, new_n_n532_, new_nt32_,
    new_nd33_, new_n_n505_, new_n_n498_, new_n_n491_, new_ne34_, new_nh34_,
    new_nr34_, new_n_n478_, new_ne35_, new_n_n453_, new_n_n444_,
    new_n_n435_, new_n_n424_, new_n_n421_, new_n_n410_, new_n_n400_,
    new_n_n389_, new_n_n360_, new_n_n349_, new_n_n338_, new_n_n327_,
    new_n_n324_, new_n_n313_, new_n_n302_, new_n_n291_, new_n_n275_,
    new_n_n261_, new_n_n250_, new_n_n239_, new_n_n228_, new_n_n214_,
    new_n_n203_, new_n_n192_, new_n_n176_, new_n_n165_, new_n_n162_,
    new_n_n151_, new_n_n140_, new_n_n129_, new_n_n104_, new_n_n93_,
    new_n_n1_, new_n_n1104_, new_n_n1064_, new_n_n1043_, new_n_n1036_,
    new_n_n1025_, new_n_n1017_, new_n_n990_, new_n_n982_, new_n_n970_,
    new_n_n962_, new_n_n958_, new_n_n950_, new_n_n938_, new_n_n930_,
    new_n_n907_, new_n_n903_, new_n_n895_, new_n_n883_, new_n_n875_,
    new_no7_, new_n_n851_, new_n_n843_, new_n_n828_, new_nz7_, new_ne8_,
    new_n_n822_, new_no8_, new_nr8_, new_nj9_, new_n_n768_, new_nk15_,
    new_n_n732_, new_ni18_, new_n_n651_, new_nu23_, new_n_n640_,
    new_n_n634_, new_nz24_, new_no25_, new_n_n593_, new_nl26_, new_ny26_,
    new_nk28_, new_n_n580_, new_nf29_, new_nn29_, new_nr29_, new_nu29_,
    new_nc31_, new_nk31_, new_nc32_, new_n_n537_, new_n_n533_, new_nu32_,
    new_nc33_, new_nr33_, new_n_n499_, new_n_n490_, new_nd34_, new_n_n485_,
    new_nq34_, new_n_n477_, new_n_n470_, new_n_n452_, new_n_n445_,
    new_n_n434_, new_n_n425_, new_n_n420_, new_n_n411_, new_n_n399_,
    new_n_n390_, new_n_n359_, new_n_n350_, new_n_n337_, new_n_n328_,
    new_n_n323_, new_n_n314_, new_n_n301_, new_n_n292_, new_n_n265_,
    new_n_n260_, new_n_n251_, new_n_n238_, new_n_n229_, new_n_n224_,
    new_n_n202_, new_n_n193_, new_n_n175_, new_n_n166_, new_n_n161_,
    new_n_n152_, new_n_n139_, new_n_n130_, new_n_n103_, new_n_n94_,
    new_n_n2_, new_n_n1096_, new_n_n1087_, new_np6_, new_nt6_,
    new_n_n1034_, new_n_n1028_, new_n_n1018_, new_n_n989_, new_n_n979_,
    new_n_n973_, new_n_n963_, new_n_n957_, new_n_n947_, new_n_n941_,
    new_n_n931_, new_n_n918_, new_n_n908_, new_n_n902_, new_n_n892_,
    new_n_n886_, new_n_n876_, new_n_n870_, new_n_n860_, new_nr7_,
    new_n_n831_, new_ny7_, new_nf8_, new_n_n820_, new_nn8_, new_n_n808_,
    new_n_n775_, new_n_n769_, new_nt9_, new_no23_, new_nw23_, new_n_n641_,
    new_ne24_, new_n_n605_, new_np25_, new_nw25_, new_ng26_, new_nx26_,
    new_n_n575_, new_n_n568_, new_ng29_, new_n_n561_, new_no29_,
    new_n_n548_, new_nd31_, new_ns31_, new_nb32_, new_nj32_, new_np32_,
    new_n_n527_, new_nb33_, new_n_n504_, new_n_n497_, new_n_n492_,
    new_nc34_, new_n_n484_, new_nt34_, new_n_n480_, new_n_n471_, new_nk35_,
    new_n_n451_, new_n_n442_, new_n_n437_, new_n_n426_, new_n_n419_,
    new_n_n408_, new_n_n401_, new_n_n391_, new_n_n376_, new_n_n365_,
    new_n_n358_, new_n_n347_, new_n_n340_, new_n_n329_, new_n_n322_,
    new_n_n311_, new_n_n304_, new_n_n293_, new_n_n277_, new_n_n266_,
    new_n_n259_, new_n_n248_, new_n_n241_, new_n_n230_, new_n_n223_,
    new_n_n212_, new_n_n194_, new_n_n178_, new_n_n167_, new_n_n160_,
    new_n_n149_, new_n_n142_, new_n_n131_, new_n_n124_, new_n_n113_,
    new_n_n3_, new_n_n1095_, new_n_n1088_, new_n_n1049_, new_n_n1042_,
    new_nv6_, new_n_n1027_, new_n_n1019_, new_n_n988_, new_n_n980_,
    new_n_n972_, new_n_n964_, new_n_n956_, new_n_n948_, new_n_n940_,
    new_n_n932_, new_n_n917_, new_n_n909_, new_n_n901_, new_n_n893_,
    new_n_n885_, new_n_n877_, new_n_n869_, new_n_n861_, new_nq7_,
    new_n_n830_, new_nx7_, new_ng8_, new_n_n821_, new_n_n815_, new_n_n809_,
    new_ni9_, new_nm9_, new_n_n764_, new_np23_, new_n_n647_, new_nz23_,
    new_nd24_, new_nj25_, new_nq25_, new_nt25_, new_ni26_, new_nv26_,
    new_n_n574_, new_na29_, new_ni29_, new_n_n562_, new_np29_, new_n_n549_,
    new_nm31_, new_nt31_, new_n_n538_, new_nk32_, new_no32_, new_ns32_,
    new_na33_, new_n_n503_, new_nv33_, new_ny33_, new_nb34_, new_ni34_,
    new_ns34_, new_n_n479_, new_nd35_, new_n_n459_, new_n_n450_,
    new_n_n443_, new_n_n436_, new_n_n427_, new_n_n418_, new_n_n409_,
    new_nh6_, new_n_n392_, new_n_n375_, new_n_n366_, new_n_n357_,
    new_n_n348_, new_n_n339_, new_n_n330_, new_n_n321_, new_n_n312_,
    new_n_n303_, new_n_n294_, new_n_n276_, new_n_n267_, new_n_n258_,
    new_n_n249_, new_n_n240_, new_n_n231_, new_n_n222_, new_n_n213_,
    new_n_n204_, new_n_n177_, new_n_n168_, new_n_n159_, new_n_n150_,
    new_n_n141_, new_n_n132_, new_n_n123_, new_n_n114_, new_n_n4_,
    new_n_n1097_, new_nv4_, new_nq6_, new_n_n1048_, new_n_n1038_,
    new_n_n1030_, new_n_n1020_, new_ng7_, new_n_n933_, new_n_n79_,
    new_n_n68_, new_n_n57_, new_n_n46_, new_n_n35_, new_nr4_, new_n_n1089_,
    new_n_n1063_, new_n_n1047_, new_n_n1039_, new_n_n1029_, new_n_n1021_,
    new_n_n942_, new_nh7_, new_n_n80_, new_n_n67_, new_n_n58_, new_n_n45_,
    new_n_n36_, new_np4_, new_n_n1099_, new_n_n1090_, new_ne5_,
    new_n_n1046_, new_nu6_, new_n_n1032_, new_n_n1022_, new_ne7_,
    new_n_n951_, new_n_n81_, new_n_n66_, new_n_n55_, new_n_n48_,
    new_n_n37_, new_n_n1098_, new_n_n1091_, new_n_n1071_, new_n_n1045_,
    new_n_n1037_, new_n_n1031_, new_n_n1023_, new_n_n960_, new_nf7_,
    new_n_n82_, new_n_n65_, new_n_n56_, new_n_n47_, new_n_n38_, new_n_n0_,
    new_nq4_, new_n_n1092_, new_nb5_, new_ng5_, new_n_n1060_, new_n_n1054_,
    new_nx6_, new_nc7_, new_n_n969_, new_nh18_, new_n_n725_, new_n_n646_,
    new_nc24_, new_no26_, new_n_n83_, new_n_n28_, new_nc6_, new_no5_,
    new_n_n10_, new_n_n1100_, new_ns4_, new_n_n1070_, new_nf5_,
    new_n_n1059_, new_nr6_, new_nw6_, new_n_n978_, new_nd7_, new_n_n729_,
    new_nr18_, new_n_n645_, new_n_n639_, new_nz25_, new_n_n84_, new_n_n27_,
    new_nd6_, new_nn5_, new_n_n11_, new_n_n1102_, new_n_n1093_,
    new_n_n1069_, new_ni5_, new_n_n1062_, new_n_n1055_, new_n_n1040_,
    new_na7_, new_n_n987_, new_n_n771_, new_n_n730_, new_np18_, new_nj23_,
    new_n_n650_, new_n_n597_, new_n_n26_, new_na6_, new_nq5_, new_n_n12_,
    new_n_n1101_, new_n_n1094_, new_n_n1068_, new_nh5_, new_n_n1061_,
    new_n_n1056_, new_ns6_, new_n_n996_, new_nb7_, new_n_n765_, new_nf18_,
    new_n_n726_, new_n_n656_, new_nq23_, new_nk25_, new_n_n25_, new_nb6_,
    new_np5_, new_n_n13_, new_n_n1084_, new_n_n1076_, new_ny6_,
    new_n_n1005_, new_n_n758_, new_n_n722_, new_nj19_, new_nv19_,
    new_n_n709_, new_n_n667_, new_nc23_, new_n_n604_, new_n_n54_,
    new_n_n43_, new_n_n32_, new_ng6_, new_n_n20_, new_n_n14_, new_n_n1083_,
    new_nz4_, new_n_n1014_, new_nz6_, new_nj15_, new_nz18_, new_n_n718_,
    new_n_n713_, new_nf20_, new_nu22_, new_nb23_, new_nw16_, new_n_n53_,
    new_n_n44_, new_n_n31_, new_n_n22_, new_nr5_, new_n_n15_, new_nw4_,
    new_n_n1077_, new_nx15_, new_nb19_, new_n_n717_, new_n_n714_,
    new_nd20_, new_n_n679_, new_n_n672_, new_n_n612_, new_n_n74_,
    new_n_n63_, new_n_n30_, new_ne6_, new_nx5_, new_n_n16_, new_n_n1085_,
    new_n_n1078_, new_n_n747_, new_n_n721_, new_nl19_, new_nt19_,
    new_n_n710_, new_n_n678_, new_n_n673_, new_n_n619_, new_n_n73_,
    new_n_n64_, new_n_n29_, new_nf6_, new_n_n21_, new_n_n17_, new_n_n1079_,
    new_ns16_, new_n_n706_, new_nx20_, new_nh21_, new_n_n691_, new_n_n690_,
    new_n_n684_, new_n_n626_, new_n_n75_, new_n_n72_, new_n_n61_,
    new_n_n50_, new_n_n39_, new_nz5_, new_n_n18_, new_n_n1086_,
    new_n_n741_, new_nn20_, new_n_n702_, new_n_n696_, new_nq21_, new_nr21_,
    new_ny21_, new_ng24_, new_n_n76_, new_n_n71_, new_n_n62_, new_n_n49_,
    new_n_n40_, new_ny5_, new_n_n19_, new_n_n737_, new_np20_, new_n_n701_,
    new_n_n698_, new_nl21_, new_n_n77_, new_n_n70_, new_n_n59_, new_n_n52_,
    new_n_n41_, new_n_n34_, new_n_n23_, new_n_n733_, new_n_n705_,
    new_nz20_, new_n_n697_, new_nk21_, new_n_n78_, new_n_n69_, new_n_n60_,
    new_n_n51_, new_n_n42_, new_n_n33_, new_n_n24_;
  assign new_na1_ = pa1;
  assign new_nb2_ = pb2;
  assign new_nc3_ = pc3;
  assign new_nd4_ = pd4;
  assign pe5 = new_ne5_;
  assign pf6 = new_nf6_;
  assign pg7 = new_ng7_;
  assign ph8 = new_nh8_;
  assign pi9 = new_ni9_;
  assign new_np_ = pp;
  assign new_na0_ = pa0;
  assign new_nb3_ = pb3;
  assign new_nc2_ = pc2;
  assign pd5 = new_nd5_;
  assign new_ne4_ = pe4;
  assign pf7 = new_nf7_;
  assign pg6 = new_ng6_;
  assign ph9 = new_nh9_;
  assign pi8 = new_ni8_;
  assign new_nq_ = pq;
  assign new_na3_ = pa3;
  assign new_nb0_ = pb0;
  assign new_nc1_ = pc1;
  assign pd6 = new_nd6_;
  assign pe7 = new_ne7_;
  assign new_nf4_ = pf4;
  assign pg5 = new_ng5_;
  assign pj8 = new_nj8_;
  assign pk9 = new_nk9_;
  assign new_nr_ = pr;
  assign new_na2_ = pa2;
  assign new_nb1_ = pb1;
  assign new_nc0_ = pc0;
  assign pd7 = new_nd7_;
  assign pe6 = new_ne6_;
  assign pf5 = new_nf5_;
  assign new_ng4_ = pg4;
  assign pj9 = new_nj9_;
  assign pk8 = new_nk8_;
  assign new_ns_ = ps;
  assign pa5 = new_na5_;
  assign pb6 = new_nb6_;
  assign pc7 = new_nc7_;
  assign new_nd0_ = pd0;
  assign new_ne1_ = pe1;
  assign new_nf2_ = pf2;
  assign new_ng3_ = pg3;
  assign pl8 = new_nl8_;
  assign pm9 = new_nm9_;
  assign new_nt_ = pt;
  assign new_na4_ = pa4;
  assign pb7 = new_nb7_;
  assign pc6 = new_nc6_;
  assign new_nd1_ = pd1;
  assign new_ne0_ = pe0;
  assign new_nf3_ = pf3;
  assign new_ng2_ = pg2;
  assign pl9 = new_nl9_;
  assign pm8 = new_nm8_;
  assign new_nu_ = pu;
  assign pa7 = new_na7_;
  assign new_nb4_ = pb4;
  assign pc5 = new_nc5_;
  assign new_nd2_ = pd2;
  assign new_ne3_ = pe3;
  assign new_nf0_ = pf0;
  assign new_ng1_ = pg1;
  assign pn8 = new_nn8_;
  assign po9 = new_no9_;
  assign new_nv_ = pv;
  assign pa6 = new_na6_;
  assign pb5 = new_nb5_;
  assign new_nc4_ = pc4;
  assign new_nd3_ = pd3;
  assign new_ne2_ = pe2;
  assign new_nf1_ = pf1;
  assign new_ng0_ = pg0;
  assign pn9 = new_nn9_;
  assign po8 = new_no8_;
  assign new_nw_ = pw;
  assign pa9 = new_na9_;
  assign new_nh0_ = ph0;
  assign new_ni1_ = pi1;
  assign new_nj2_ = pj2;
  assign new_nk3_ = pk3;
  assign new_nl4_ = pl4;
  assign pm5 = new_nm4_;
  assign pn6 = new_nn6_;
  assign po7 = new_no7_;
  assign new_nx_ = px;
  assign pa8 = new_na8_;
  assign new_nh1_ = ph1;
  assign new_ni0_ = pi0;
  assign new_nj3_ = pj3;
  assign new_nk2_ = pk2;
  assign pl5 = new_nl5_;
  assign new_nm4_ = pm4;
  assign pn7 = new_nn7_;
  assign po6 = new_no6_;
  assign new_ny_ = py;
  assign pb8 = new_nb8_;
  assign pc9 = new_nc9_;
  assign new_nh2_ = ph2;
  assign new_ni3_ = pi3;
  assign new_nj0_ = pj0;
  assign new_nk1_ = pk1;
  assign pl6 = new_nl6_;
  assign pm7 = new_nm7_;
  assign new_nn4_ = pn4;
  assign po5 = new_no5_;
  assign new_nz_ = pz;
  assign pb9 = new_nb9_;
  assign pc8 = new_nc8_;
  assign new_nh3_ = ph3;
  assign new_ni2_ = pi2;
  assign new_nj1_ = pj1;
  assign new_nk0_ = pk0;
  assign pl7 = new_nl7_;
  assign pm6 = new_nk4_;
  assign pn5 = new_nn5_;
  assign po4 = new_no4_;
  assign pd8 = new_nd8_;
  assign pe9 = new_ne9_;
  assign new_nh4_ = ph4;
  assign pi5 = new_ni5_;
  assign pj6 = new_nj6_;
  assign pk7 = new_nk7_;
  assign new_nl0_ = pl0;
  assign new_nm1_ = pm1;
  assign new_nn2_ = pn2;
  assign new_no3_ = po3;
  assign pd9 = new_nd9_;
  assign pe8 = new_ne8_;
  assign ph5 = new_nh5_;
  assign new_ni4_ = pi4;
  assign pj7 = new_nj7_;
  assign pk6 = new_nk6_;
  assign new_nl1_ = pl1;
  assign new_nm0_ = pm0;
  assign new_nn3_ = pn3;
  assign new_no2_ = po2;
  assign pf8 = new_nf8_;
  assign pg9 = new_ng9_;
  assign ph6 = new_nh6_;
  assign pi7 = new_ni7_;
  assign new_nj4_ = pj4;
  assign pk5 = new_nk5_;
  assign new_nl2_ = pl2;
  assign new_nm3_ = pm3;
  assign new_nn0_ = pn0;
  assign new_no1_ = po1;
  assign pf9 = new_nf9_;
  assign pg8 = new_ng8_;
  assign ph7 = new_nh7_;
  assign pi6 = new_ni6_;
  assign pj5 = new_nj5_;
  assign new_nk4_ = pk4;
  assign new_nl3_ = pl3;
  assign new_nm2_ = pm2;
  assign new_nn1_ = pn1;
  assign new_no0_ = po0;
  assign new_np0_ = pp0;
  assign new_nq1_ = pq1;
  assign new_nr2_ = pr2;
  assign new_ns3_ = ps3;
  assign pt4 = new_nu3_;
  assign pu5 = new_nw5_;
  assign pv6 = new_nv6_;
  assign pw7 = new_nw7_;
  assign px8 = new_nx8_;
  assign new_na_ = pa;
  assign new_np1_ = pp1;
  assign new_nq0_ = pq0;
  assign new_nr3_ = pr3;
  assign new_ns2_ = ps2;
  assign pt5 = new_nw5_;
  assign pu4 = new_nv3_;
  assign pv7 = new_nv7_;
  assign pw6 = new_nw6_;
  assign py8 = new_ny8_;
  assign new_nb_ = pb;
  assign new_np2_ = pp2;
  assign new_nq3_ = pq3;
  assign new_ns1_ = ps1;
  assign pt6 = new_nt6_;
  assign pu7 = new_nu7_;
  assign pv4 = new_nv4_;
  assign pw5 = new_nw5_;
  assign pz8 = new_nz8_;
  assign new_nc_ = pc;
  assign new_np3_ = pp3;
  assign new_nq2_ = pq2;
  assign new_nr1_ = pr1;
  assign new_ns0_ = ps0;
  assign pt7 = new_nt7_;
  assign pu6 = new_nu6_;
  assign pv5 = new_nw5_;
  assign pw4 = new_nw4_;
  assign new_nd_ = pd;
  assign pp4 = new_np4_;
  assign pq5 = new_nq5_;
  assign pr6 = new_nr6_;
  assign ps7 = new_ns7_;
  assign new_nt0_ = pt0;
  assign new_nu1_ = pu1;
  assign new_nv2_ = pv2;
  assign new_nw3_ = pw3;
  assign new_ne_ = pe;
  assign pp5 = new_np5_;
  assign pq4 = new_nq4_;
  assign pr7 = new_nr7_;
  assign ps6 = new_ns6_;
  assign new_nt1_ = pt1;
  assign new_nu0_ = pu0;
  assign new_nv3_ = pv3;
  assign new_nw2_ = pw2;
  assign new_nf_ = pf;
  assign pp6 = new_np6_;
  assign pq7 = new_nq7_;
  assign pr4 = new_nr4_;
  assign ps5 = new_nw5_;
  assign new_nt2_ = pt2;
  assign new_nu3_ = pu3;
  assign new_nv0_ = pv0;
  assign new_nw1_ = pw1;
  assign new_ng_ = pg;
  assign pp7 = new_np7_;
  assign pq6 = new_nq6_;
  assign pr5 = new_nr5_;
  assign ps4 = new_ns4_;
  assign new_nt3_ = pt3;
  assign new_nu2_ = pu2;
  assign new_nv1_ = pv1;
  assign new_nw0_ = pw0;
  assign new_nh_ = ph;
  assign pp8 = new_np8_;
  assign pq9 = new_nq9_;
  assign new_nx0_ = px0;
  assign new_ny1_ = py1;
  assign new_nz2_ = pz2;
  assign new_ni_ = pi;
  assign pp9 = new_np9_;
  assign pq8 = new_nq8_;
  assign new_nx1_ = px1;
  assign new_ny0_ = py0;
  assign new_nz3_ = pz3;
  assign new_nj_ = pj;
  assign pr8 = new_nr8_;
  assign ps9 = new_ns9_;
  assign new_nx2_ = px2;
  assign new_ny3_ = py3;
  assign new_nz0_ = pz0;
  assign new_nk_ = pk;
  assign pr9 = new_nr9_;
  assign ps8 = new_ns8_;
  assign new_nx3_ = px3;
  assign new_ny2_ = py2;
  assign new_nz1_ = pz1;
  assign new_nl_ = pl;
  assign pt8 = new_nt8_;
  assign pu9 = new_nu9_;
  assign px4 = new_nx4_;
  assign py5 = new_ny5_;
  assign pz6 = new_nz6_;
  assign new_nm_ = pm;
  assign pt9 = new_nt9_;
  assign pu8 = new_nu8_;
  assign px5 = new_nx5_;
  assign py4 = new_ny4_;
  assign pz7 = new_nz7_;
  assign new_nn_ = pn;
  assign pv8 = new_nv8_;
  assign pw9 = new_nw9_;
  assign px6 = new_nx6_;
  assign py7 = new_ny7_;
  assign pz4 = new_nz4_;
  assign new_no_ = po;
  assign pv9 = new_nv9_;
  assign pw8 = new_nw8_;
  assign px7 = new_nx7_;
  assign py6 = new_ny6_;
  assign pz5 = new_nz5_;
  assign new_n_n1007_ = new_n_n41_ & new_n_n83_ & new_n_n42_;
  assign new_n_n997_ = new_n_n350_ & new_n_n83_ & new_n_n44_;
  assign new_n_n920_ = new_n_n61_ & new_n_n432_ & new_n_n62_;
  assign new_n_n910_ = new_n_n350_ & new_n_n432_ & new_n_n64_;
  assign new_n_n900_ = new_na17_ & new_n_n83_ & new_n_n66_;
  assign new_n_n890_ = new_n_n67_ & new_n_n83_ & new_n_n68_;
  assign new_n_n880_ = new_n_n350_ & new_n_n83_ & new_n_n70_;
  assign new_n_n833_ = new_n_n81_ & new_nj2_ & new_n_n82_;
  assign new_nw7_ = new_n_n408_ & new_no0_ & new_n_n87_;
  assign new_nh8_ = new_n_n408_ & new_no0_ & new_n_n98_;
  assign new_n_n819_ = new_n_n194_ & new_n_n107_ & new_n_n145_;
  assign new_np8_ = new_n_n810_ | new_n_n811_;
  assign new_n_n804_ = new_no0_ & new_n_n122_ & new_n_n147_;
  assign new_n_n797_ = new_n_n194_ & new_n_n129_ & new_n_n145_;
  assign new_na9_ = new_n_n788_ | new_n_n789_;
  assign new_n_n770_ = new_no0_ & new_n_n166_ & new_n_n165_;
  assign new_nq9_ = new_n_n179_ | new_n_n763_ | new_n_n762_;
  assign new_nv9_ = new_n_n756_ | new_n_n757_;
  assign new_no15_ = new_n_n752_ | new_n_n753_;
  assign new_n_n749_ = new_n_n204_ & new_nc1_;
  assign new_nm16_ = new_n_n205_ & new_nt15_;
  assign new_na17_ = new_n_n434_ & new_n_n433_ & new_n_n209_;
  assign new_nl17_ = new_n_n217_ & new_nl4_;
  assign new_nx17_ = new_n_n733_ | new_n_n218_;
  assign new_nm19_ = new_n_n716_ | new_n_n742_ | new_n_n697_;
  assign new_n_n712_ = new_nv_ & new_no0_ & new_n_n408_;
  assign new_ni20_ = new_n_n247_ & new_nl4_;
  assign new_nu20_ = new_n_n703_ | new_n_n248_;
  assign new_n_n699_ = new_n_n255_ & new_n_n378_ & new_n_n254_;
  assign new_nj21_ = new_nl2_ | new_n_n365_;
  assign new_n_n687_ = new_nk0_ & new_n_n430_ & new_nj_;
  assign new_na22_ = new_nm2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n676_ = new_n_n428_ & new_n_n350_ & new_n_n269_;
  assign new_nt22_ = new_n_n669_ | new_n_n668_ | new_n_n667_;
  assign new_n_n663_ = new_ng_ & new_nl0_;
  assign new_ni23_ = new_ns2_ | new_n_n365_;
  assign new_n_n630_ = new_n_n292_ & new_n_n294_ & new_n_n293_;
  assign new_nl24_ = new_nx2_ & new_nl4_;
  assign new_n_n616_ = new_nn_ & new_n_n305_ & new_n_n353_;
  assign new_nw24_ = new_nn0_ | new_nm0_ | new_n_n307_;
  assign new_nd25_ = new_nq0_ | new_n_n419_;
  assign new_n_n600_ = new_nj6_ & new_n_n404_ & new_n_n313_;
  assign new_nr25_ = new_n_n597_ | new_n_n596_ | new_n_n595_;
  assign new_ng27_ = new_n_n439_ | new_n_n322_ | new_nj25_;
  assign new_nw27_ = new_nq0_ | new_n_n416_;
  assign new_n_n590_ = new_nh1_ & new_n_n326_;
  assign new_nm28_ = new_n_n439_ | new_nj25_ | new_n_n331_;
  assign new_nu28_ = new_n_n571_ | new_n_n570_ | new_n_n576_ | new_n_n569_ | new_n_n573_ | new_n_n572_ | new_n_n575_ | new_n_n574_;
  assign new_nx28_ = new_nk6_ | new_nj1_ | new_n_n394_;
  assign new_nj29_ = new_n_n564_ | new_n_n565_;
  assign new_n_n559_ = new_n_n347_ & new_n_n432_ & new_n_n348_;
  assign new_na30_ = new_nq0_ | new_n_n433_;
  assign new_nl30_ = new_n_n546_ | new_nz29_;
  assign new_n_n544_ = new_n_n404_ & new_nl25_ & new_n_n367_;
  assign new_ni31_ = new_n_n408_ & new_no4_ & new_n_n372_;
  assign new_n_n541_ = new_nl25_ & new_n_n377_ & new_n_n376_;
  assign new_na32_ = new_n_n538_ | new_nz29_;
  assign new_nl32_ = new_ng1_ | new_nj25_ | new_n_n412_;
  assign new_n_n530_ = new_nl6_ & new_n_n394_;
  assign new_nx32_ = new_n_n524_ | new_n_n525_;
  assign new_nh33_ = new_n_n521_ | new_n_n520_ | new_n_n517_;
  assign new_nl33_ = new_n_n514_ | new_n_n513_ | new_n_n512_;
  assign new_n_n507_ = new_n_n426_ & new_n_n417_;
  assign new_n_n501_ = new_nk0_ & new_nl0_ & new_n_n421_;
  assign new_nx33_ = new_n_n428_ | new_n_n493_ | new_n_n492_;
  assign new_n_n486_ = new_n_n431_ & new_n_n430_ & new_n_n429_;
  assign new_nk34_ = new_n_n439_ & new_nm1_ & new_nh1_;
  assign new_nw34_ = new_nz3_ & new_n_n441_;
  assign new_n_n475_ = new_ni6_ & new_nj6_ & new_n_n442_;
  assign new_n_n469_ = new_n_n447_ & new_n_n450_;
  assign new_nl35_ = new_n_n454_ | new_ng1_ | new_n_n455_;
  assign new_n_n457_ = ~new_nh4_;
  assign new_nj6_ = ~new_nj1_;
  assign new_n_n439_ = ~new_nk4_;
  assign new_n_n428_ = ~new_nm0_;
  assign new_n_n417_ = ~new_nb3_;
  assign new_n_n406_ = ~new_nb33_;
  assign new_n_n396_ = ~new_nq25_;
  assign new_no4_ = ~new_ng1_;
  assign new_n_n364_ = ~new_nn30_;
  assign new_n_n353_ = ~new_ns23_;
  assign new_n_n342_ = ~new_ng29_;
  assign new_n_n331_ = ~new_nn28_;
  assign new_n_n320_ = ~new_nm3_;
  assign new_n_n309_ = ~new_nr25_;
  assign new_n_n298_ = ~new_nx2_;
  assign new_n_n287_ = ~new_na24_;
  assign new_n_n254_ = ~new_nw16_;
  assign new_n_n243_ = ~new_ne2_;
  assign new_n_n232_ = ~new_nh19_;
  assign new_n_n221_ = ~new_nt1_;
  assign new_n_n210_ = ~new_ne17_;
  assign new_n_n199_ = ~new_nz15_;
  assign new_n_n188_ = ~new_nn32_;
  assign new_n_n144_ = ~new_nc28_;
  assign new_n_n133_ = ~new_nm27_;
  assign new_n_n122_ = ~new_nv26_;
  assign new_n_n111_ = ~new_nf26_;
  assign new_n_n100_ = ~new_nw24_;
  assign new_n_n89_ = ~new_ns22_;
  assign new_n_n1006_ = new_n_n350_ & new_n_n83_ & new_n_n42_;
  assign new_n_n998_ = new_n_n43_ & new_n_n83_ & new_n_n44_;
  assign new_n_n919_ = new_n_n350_ & new_n_n432_ & new_n_n62_;
  assign new_n_n911_ = new_n_n63_ & new_n_n432_ & new_n_n64_;
  assign new_n_n899_ = new_n_n65_ & new_n_n83_ & new_n_n66_;
  assign new_n_n891_ = new_na17_ & new_n_n83_ & new_n_n68_;
  assign new_n_n871_ = new_n_n350_ & new_n_n83_ & new_n_n72_;
  assign new_n_n832_ = new_n_n350_ & new_nj2_ & new_n_n82_;
  assign new_nv7_ = new_n_n408_ & new_no0_ & new_n_n86_;
  assign new_ni8_ = new_n_n824_ | new_n_n825_;
  assign new_nl8_ = new_n_n818_ | new_n_n819_;
  assign new_n_n811_ = new_n_n194_ & new_n_n115_ & new_n_n145_;
  assign new_n_n805_ = new_n_n194_ & new_n_n121_ & new_n_n145_;
  assign new_n_n796_ = new_no0_ & new_n_n130_ & new_n_n147_;
  assign new_n_n790_ = new_no0_ & new_n_n136_ & new_n_n147_;
  assign new_nh9_ = new_n_n411_ | new_n_n154_ | new_n_n775_;
  assign new_n_n763_ = new_n_n181_ & new_n_n194_ & new_n_n180_;
  assign new_nu9_ = new_n_n191_ & new_nm1_;
  assign new_n_n753_ = new_ne1_ & new_nd1_;
  assign new_n_n750_ = new_n_n205_ & new_n_n201_;
  assign new_np16_ = new_nq0_ | new_n_n411_ | new_n_n745_;
  assign new_n_n742_ = new_nn0_ & new_no0_ & new_n_n408_;
  assign new_nn17_ = new_n_n737_ | new_n_n214_;
  assign new_nv17_ = new_n_n221_ & new_nl4_;
  assign new_n_n716_ = new_nt_ & new_no0_ & new_n_n408_;
  assign new_nw19_ = new_n_n712_ | new_n_n742_ | new_n_n697_;
  assign new_nk20_ = new_n_n707_ | new_n_n244_;
  assign new_ns20_ = new_n_n251_ & new_nl4_;
  assign new_nf21_ = new_n_n698_ | new_n_n742_ | new_n_n697_;
  assign new_n_n692_ = new_nk0_ & new_n_n430_ & new_ni_;
  assign new_ns21_ = new_nm2_ | new_n_n365_;
  assign new_nz21_ = new_nn2_ | new_n_n365_;
  assign new_n_n675_ = new_n_n387_ & new_n_n270_ & new_n_n279_;
  assign new_n_n670_ = new_n_n387_ & new_n_n273_ & new_n_n279_;
  assign new_n_n662_ = new_nk0_ & new_n_n430_ & new_no_;
  assign new_n_n657_ = new_nk0_ & new_n_n430_ & new_np_;
  assign new_n_n629_ = new_n_n387_ & new_n_n294_ & new_n_n293_;
  assign new_n_n623_ = new_n_n387_ & new_n_n297_ & new_n_n296_;
  assign new_n_n615_ = new_n_n365_ & new_nx2_ & new_n_n306_;
  assign new_n_n609_ = new_n_n365_ & new_ny2_ & new_n_n306_;
  assign new_ne25_ = new_n_n602_ | new_n_n604_ | new_n_n603_ | new_n_n605_;
  assign new_n_n601_ = new_nl6_ & new_n_n404_ & new_n_n313_;
  assign new_nx25_ = new_nq0_ | new_n_n417_;
  assign new_nh27_ = new_nq0_ | new_n_n321_;
  assign new_nv27_ = new_n_n439_ | new_n_n414_ | new_nj25_;
  assign new_n_n589_ = new_nh1_ & new_n_n396_;
  assign new_n_n582_ = new_n_n330_ & new_n_n335_ & new_n_n329_;
  assign new_n_n576_ = new_n_n400_ & new_n_n393_ & new_n_n336_;
  assign new_nw28_ = new_n_n339_ & new_nl6_;
  assign new_n_n565_ = new_n_n378_ & new_n_n408_ & new_n_n344_;
  assign new_n_n560_ = new_n_n346_ & new_n_n432_ & new_n_n348_;
  assign new_nb30_ = new_n_n547_ | new_nz29_;
  assign new_nk30_ = new_nq0_ | new_n_n434_;
  assign new_nv30_ = new_nq0_ | new_n_n378_;
  assign new_nh31_ = new_n_n404_ & new_nl25_ & new_n_n371_;
  assign new_nr31_ = new_n_n378_ | new_nq0_ | new_n_n379_;
  assign new_nz31_ = new_n_n457_ | new_ng1_ | new_nq0_;
  assign new_nm32_ = new_n_n405_ | new_ng1_ | new_nq0_;
  assign new_n_n531_ = new_nk6_ & new_n_n393_;
  assign new_n_n522_ = new_nd33_ & new_n_n412_;
  assign new_n_n521_ = new_n_n413_ & new_n_n430_;
  assign new_n_n515_ = new_n_n427_ & new_nl0_;
  assign new_np33_ = new_n_n428_ & new_n_n418_;
  assign new_nt33_ = new_n_n428_ | new_n_n501_ | new_n_n500_;
  assign new_n_n493_ = new_nk0_ & new_nl0_ & new_n_n425_;
  assign new_n_n487_ = new_nk0_ & new_nl0_ & new_n_n429_;
  assign new_nl34_ = new_n_n439_ & new_nm1_ & new_ni1_;
  assign new_nv34_ = new_n_n458_ | new_n_n440_ | new_n_n459_;
  assign new_n_n474_ = new_ny0_ & new_nj6_ & new_n_n442_;
  assign new_nh35_ = new_n_n468_ | new_n_n466_ | new_n_n465_ | new_n_n467_ | new_n_n469_;
  assign new_n_n468_ = new_nj6_ & new_nk6_ & new_n_n447_;
  assign new_n_n456_ = ~new_ng4_;
  assign new_n_n447_ = ~new_nj35_;
  assign new_n_n438_ = ~new_ng34_;
  assign new_n_n429_ = ~new_nl3_;
  assign new_n_n416_ = ~new_ns3_;
  assign new_n_n407_ = ~new_nq30_;
  assign new_n_n395_ = ~new_ns0_;
  assign new_n_n386_ = ~new_nj32_;
  assign new_n_n363_ = ~new_no30_;
  assign new_n_n354_ = ~new_nv29_;
  assign new_n_n341_ = ~new_nf29_;
  assign new_n_n332_ = ~new_np28_;
  assign new_n_n319_ = ~new_ns25_;
  assign new_n_n310_ = ~new_np25_;
  assign new_n_n297_ = ~new_nl24_;
  assign new_n_n288_ = ~new_nz23_;
  assign new_n_n264_ = ~new_nz21_;
  assign new_n_n242_ = ~new_ng20_;
  assign new_n_n233_ = ~new_nz1_;
  assign new_n_n220_ = ~new_nd18_;
  assign new_n_n211_ = ~new_no1_;
  assign new_n_n198_ = ~new_np35_;
  assign new_n_n189_ = ~new_nm32_;
  assign new_n_n143_ = ~new_nb28_;
  assign new_n_n134_ = ~new_nn27_;
  assign new_n_n121_ = ~new_nu26_;
  assign new_n_n112_ = ~new_ng26_;
  assign new_n_n99_ = ~new_nx24_;
  assign new_n_n90_ = ~new_nz22_;
  assign new_ny4_ = new_n_n1079_ | new_n_n1078_ | new_n_n1077_;
  assign new_n_n1009_ = new_n_n350_ & new_n_n432_ & new_n_n42_;
  assign new_n_n999_ = new_na17_ & new_n_n83_ & new_n_n44_;
  assign new_n_n922_ = new_n_n350_ & new_nz1_ & new_n_n62_;
  assign new_n_n912_ = new_na17_ & new_n_n432_ & new_n_n64_;
  assign new_n_n898_ = new_n_n350_ & new_n_n83_ & new_n_n66_;
  assign new_n_n882_ = new_na17_ & new_n_n83_ & new_n_n70_;
  assign new_n_n872_ = new_n_n71_ & new_n_n83_ & new_n_n72_;
  assign new_ns7_ = new_n_n833_ | new_n_n831_ | new_n_n830_ | new_n_n832_ | new_n_n834_ | new_n_n829_ | new_n_n828_ | new_n_n827_ | new_n_n826_;
  assign new_nu7_ = new_n_n408_ & new_no0_ & new_n_n85_;
  assign new_n_n825_ = new_n_n100_ & new_n_n99_ & new_n_n353_;
  assign new_nm8_ = new_n_n816_ | new_n_n817_;
  assign new_n_n813_ = new_n_n194_ & new_n_n113_ & new_n_n145_;
  assign new_ns8_ = new_n_n804_ | new_n_n805_;
  assign new_nd9_ = new_n_n782_ | new_n_n783_;
  assign new_n_n776_ = new_nl4_ & new_n_n387_ & new_n_n153_;
  assign new_n_n762_ = new_no0_ & new_n_n183_ & new_n_n182_;
  assign new_n_n756_ = new_n_n192_ & new_n_n193_;
  assign new_nl15_ = new_nh6_ | new_ng1_ | new_nq0_;
  assign new_nb16_ = new_n_n750_ | new_n_n749_ | new_n_n747_;
  assign new_n_n745_ = new_nm1_ & new_n_n206_;
  assign new_nd17_ = new_n_n741_ | new_n_n210_;
  assign new_nj17_ = new_n_n738_ | new_n_n742_ | new_n_n697_;
  assign new_n_n734_ = new_nf0_ & new_no0_ & new_n_n408_;
  assign new_ns18_ = new_n_n724_ | new_n_n742_ | new_n_n697_;
  assign new_n_n720_ = new_nr_ & new_no0_ & new_n_n408_;
  assign new_n_n707_ = new_n_n245_ & new_n_n378_ & new_n_n254_;
  assign new_nv20_ = new_n_n702_ | new_n_n742_ | new_n_n697_;
  assign new_nc21_ = new_n_n252_ & new_nl4_;
  assign new_n_n693_ = new_na_ & new_nl0_;
  assign new_n_n689_ = new_nb_ & new_n_n431_;
  assign new_n_n682_ = new_nk0_ & new_n_n430_ & new_nk_;
  assign new_nm22_ = new_n_n674_ | new_n_n673_ | new_n_n672_;
  assign new_n_n668_ = new_nf_ & new_nl0_;
  assign new_na23_ = new_n_n664_ | new_n_n663_ | new_n_n662_;
  assign new_n_n658_ = new_nh_ & new_nl0_;
  assign new_n_n632_ = new_n_n293_ & new_n_n301_;
  assign new_n_n624_ = new_n_n295_ & new_n_n297_ & new_n_n296_;
  assign new_ns24_ = new_n_n611_ | new_n_n613_ | new_n_n612_ | new_n_n614_;
  assign new_ny24_ = new_nq0_ | new_n_n308_;
  assign new_n_n607_ = new_n_n310_ & new_nh1_;
  assign new_ni25_ = new_n_n600_ | new_n_n601_;
  assign new_nm26_ = new_nq0_ | new_n_n423_;
  assign new_nd27_ = new_n_n439_ | new_n_n321_ | new_nj25_;
  assign new_nt27_ = new_nq0_ | new_n_n418_;
  assign new_n_n588_ = new_n_n327_ & new_n_n395_;
  assign new_n_n581_ = new_nl6_ & new_nl25_ & new_n_n332_;
  assign new_n_n578_ = new_n_n334_ & new_ni6_;
  assign new_nv28_ = new_nk6_ & new_nl1_;
  assign new_n_n554_ = new_nm0_ & new_na4_ & new_n_n352_;
  assign new_nx29_ = new_n_n411_ | new_n_n356_ | new_n_n357_;
  assign new_nj30_ = new_n_n411_ | new_n_n407_ | new_n_n361_;
  assign new_nw30_ = new_n_n454_ | new_n_n439_;
  assign new_n_n542_ = new_nl25_ & new_n_n377_ & new_n_n373_;
  assign new_nq31_ = new_n_n541_ | new_nz29_;
  assign new_ny31_ = new_n_n381_ | new_n_n382_ | new_n_n383_;
  assign new_nn32_ = new_n_n535_ | new_n_n533_ | new_n_n532_ | new_n_n534_ | new_n_n536_;
  assign new_nw32_ = new_n_n412_ | new_n_n403_ | new_n_n526_;
  assign new_ne33_ = new_nq0_ | new_n_n411_ | new_n_n522_;
  assign new_nq33_ = new_n_n506_ | new_n_n505_ | new_n_n502_;
  assign new_nu33_ = new_n_n428_ | new_n_n499_ | new_n_n498_;
  assign new_n_n495_ = new_nk0_ & new_nl0_ & new_n_n424_;
  assign new_na34_ = new_n_n428_ | new_n_n487_ | new_n_n486_;
  assign new_nm34_ = new_n_n439_ & new_nm1_ & new_nj1_;
  assign new_n_n483_ = new_nz0_ & new_na1_ & new_nb1_;
  assign new_n_n476_ = new_nj6_ & new_nk6_ & new_nl6_;
  assign new_ng35_ = new_nf4_ & new_ne4_ & new_n_n446_;
  assign new_n_n455_ = ~new_nm35_;
  assign new_n_n446_ = ~new_no35_;
  assign new_n_n441_ = ~new_na4_;
  assign new_n_n430_ = ~new_nl0_;
  assign new_n_n415_ = ~new_nc3_;
  assign new_n_n404_ = ~new_nj25_;
  assign new_n_n398_ = ~new_nt32_;
  assign new_n_n387_ = ~new_na17_;
  assign new_n_n362_ = ~new_np30_;
  assign new_n_n351_ = ~new_nw29_;
  assign new_n_n344_ = ~new_nk29_;
  assign new_n_n333_ = ~new_nq28_;
  assign new_n_n318_ = ~new_nn25_;
  assign new_n_n307_ = ~new_np_;
  assign new_n_n300_ = ~new_np24_;
  assign new_n_n289_ = ~new_nu2_;
  assign new_n_n263_ = ~new_ny21_;
  assign new_n_n252_ = ~new_nk2_;
  assign new_n_n234_ = ~new_nm19_;
  assign new_n_n219_ = ~new_ns1_;
  assign new_n_n208_ = ~new_nn1_;
  assign new_n_n201_ = ~new_nc1_;
  assign new_n_n190_ = ~new_na33_;
  assign new_n_n164_ = ~new_nj30_;
  assign new_n_n153_ = ~new_na29_;
  assign new_n_n120_ = ~new_ns26_;
  assign new_n_n109_ = ~new_nc26_;
  assign new_n_n102_ = ~new_ny24_;
  assign new_n_n91_ = ~new_ng23_;
  assign new_n_n1072_ = new_nk0_ & new_nl0_ & new_n_n17_;
  assign new_n_n1008_ = new_na17_ & new_n_n83_ & new_n_n42_;
  assign new_n_n1000_ = new_n_n350_ & new_n_n432_ & new_n_n44_;
  assign new_n_n921_ = new_na17_ & new_n_n432_ & new_n_n62_;
  assign new_n_n913_ = new_n_n350_ & new_na2_ & new_n_n64_;
  assign new_n_n889_ = new_n_n350_ & new_n_n83_ & new_n_n68_;
  assign new_n_n881_ = new_n_n69_ & new_n_n83_ & new_n_n70_;
  assign new_n_n873_ = new_na17_ & new_n_n83_ & new_n_n72_;
  assign new_n_n834_ = new_na17_ & new_nj2_ & new_n_n82_;
  assign new_nt7_ = new_n_n408_ & new_no0_ & new_n_n84_;
  assign new_n_n824_ = new_no0_ & new_n_n102_ & new_n_n101_;
  assign new_n_n818_ = new_no0_ & new_n_n108_ & new_n_n147_;
  assign new_n_n812_ = new_no0_ & new_n_n114_ & new_n_n147_;
  assign new_n_n806_ = new_no0_ & new_n_n120_ & new_n_n147_;
  assign new_n_n783_ = new_n_n194_ & new_n_n143_ & new_n_n145_;
  assign new_n_n777_ = new_n_n153_ & new_nx3_;
  assign new_nr9_ = new_n_n760_ | new_n_n761_;
  assign new_n_n757_ = new_n_n192_ & new_n_n206_;
  assign new_nm15_ = new_nt15_ & new_n_n432_ & new_n_n197_;
  assign new_nz15_ = new_n_n746_ | new_ni1_;
  assign new_nr16_ = new_n_n211_ & new_nl4_;
  assign new_nb17_ = new_n_n213_ & new_nl4_;
  assign new_n_n738_ = new_nh0_ & new_no0_ & new_n_n408_;
  assign new_nt17_ = new_n_n734_ | new_n_n742_ | new_n_n697_;
  assign new_n_n724_ = new_nl0_ & new_no0_ & new_n_n408_;
  assign new_nc19_ = new_n_n720_ | new_n_n742_ | new_n_n697_;
  assign new_nl20_ = new_n_n706_ | new_n_n742_ | new_n_n697_;
  assign new_n_n703_ = new_n_n249_ & new_n_n378_ & new_n_n254_;
  assign new_ne21_ = new_n_n699_ | new_n_n253_;
  assign new_n_n694_ = new_na_ & new_n_n431_;
  assign new_n_n688_ = new_nb_ & new_nl0_;
  assign new_n_n683_ = new_nc_ & new_nl0_;
  assign new_n_n674_ = new_ne_ & new_n_n431_;
  assign new_n_n669_ = new_nf_ & new_n_n431_;
  assign new_n_n664_ = new_ng_ & new_n_n431_;
  assign new_n_n659_ = new_nh_ & new_n_n431_;
  assign new_n_n631_ = new_n_n292_ & new_na17_ & new_n_n293_;
  assign new_n_n625_ = new_n_n295_ & new_na17_ & new_n_n296_;
  assign new_n_n614_ = new_n_n303_ & new_n_n301_;
  assign new_nx24_ = new_n_n378_ | new_nq0_ | new_n_n411_;
  assign new_n_n606_ = new_n_n396_ & new_ni1_;
  assign new_nh25_ = new_n_n439_ | new_n_n312_ | new_n_n526_;
  assign new_nb27_ = new_nq0_ | new_n_n429_;
  assign new_ne27_ = new_nq0_ | new_n_n320_;
  assign new_ns27_ = new_n_n439_ | new_n_n416_ | new_nj25_;
  assign new_n_n587_ = new_n_n327_ & new_n_n326_;
  assign new_nn28_ = new_n_n580_ | new_n_n581_;
  assign new_n_n577_ = new_ni1_ & new_n_n335_ & new_nt0_;
  assign new_n_n569_ = new_n_n338_ & new_n_n337_ & new_n_n336_;
  assign new_n_n553_ = new_nm0_ & new_nt15_ & new_n_n352_;
  assign new_nw29_ = new_nl4_ & new_nz3_ & new_ny3_;
  assign new_ny29_ = new_nx3_ | new_na17_ | new_nq0_;
  assign new_nx30_ = new_nk4_ & new_n_n404_ & new_nl25_;
  assign new_nj31_ = new_n_n542_ | new_nz29_;
  assign new_nz29_ = new_n_n432_ & new_nt15_;
  assign new_nw31_ = new_nk4_ & new_n_n456_ & new_nf4_;
  assign new_n_n529_ = new_nl6_ & new_nk6_;
  assign new_n_n526_ = new_nk1_ & new_nl1_;
  assign new_n_n523_ = new_n_n410_ & new_nh1_;
  assign new_n_n506_ = new_n_n419_ & new_n_n430_;
  assign new_n_n500_ = new_n_n431_ & new_n_n430_ & new_n_n421_;
  assign new_n_n494_ = new_n_n431_ & new_n_n430_ & new_n_n424_;
  assign new_n_n488_ = new_n_n431_ & new_n_n430_ & new_n_n427_;
  assign new_nn34_ = new_n_n439_ & new_nm1_ & new_nk1_;
  assign new_nx34_ = new_n_n478_ | new_n_n477_ | new_n_n483_ | new_n_n476_ | new_n_n480_ | new_n_n479_ | new_n_n482_ | new_n_n481_;
  assign new_nb35_ = new_n_n472_ | new_n_n474_ | new_n_n473_ | new_n_n475_;
  assign new_nf35_ = new_n_n456_ & new_nf4_ & new_ne4_;
  assign new_n_n454_ = ~new_nd4_;
  assign new_nk6_ = ~new_nk1_;
  assign new_n_n440_ = ~new_nx3_;
  assign new_n_n431_ = ~new_nk0_;
  assign new_n_n414_ = ~new_nt3_;
  assign new_n_n405_ = ~new_nj4_;
  assign new_n_n397_ = ~new_nu32_;
  assign new_n_n388_ = ~new_ny32_;
  assign new_n_n361_ = ~new_nr30_;
  assign new_n_n352_ = ~new_nt29_;
  assign new_n_n343_ = ~new_nm29_;
  assign new_n_n334_ = ~new_nu28_;
  assign new_n_n317_ = ~new_ny0_;
  assign new_n_n308_ = ~new_nz2_;
  assign new_n_n299_ = ~new_nq24_;
  assign new_n_n290_ = ~new_ne24_;
  assign new_n_n262_ = ~new_na22_;
  assign new_n_n253_ = ~new_nf21_;
  assign new_n_n244_ = ~new_nl20_;
  assign new_n_n218_ = ~new_ny17_;
  assign new_n_n209_ = ~new_nq35_;
  assign new_n_n200_ = ~new_nd16_;
  assign new_n_n191_ = ~new_nc33_;
  assign new_n_n163_ = ~new_ny29_;
  assign new_n_n154_ = ~new_ne29_;
  assign new_n_n119_ = ~new_nr26_;
  assign new_n_n110_ = ~new_nd26_;
  assign new_n_n101_ = ~new_nz24_;
  assign new_n_n92_ = ~new_nn23_;
  assign new_n_n1081_ = new_nk0_ & new_nl0_ & new_n_n14_;
  assign new_n_n1073_ = new_n_n17_ & new_nr3_;
  assign new_n_n1011_ = new_na17_ & new_n_n432_ & new_n_n42_;
  assign new_n_n1001_ = new_n_n43_ & new_n_n432_ & new_n_n44_;
  assign new_n_n924_ = new_na17_ & new_nz1_ & new_n_n62_;
  assign new_n_n914_ = new_n_n63_ & new_na2_ & new_n_n64_;
  assign new_n_n864_ = new_na17_ & new_n_n83_ & new_n_n74_;
  assign new_n_n854_ = new_n_n75_ & new_n_n83_ & new_n_n76_;
  assign new_n_n844_ = new_n_n350_ & new_n_n83_ & new_n_n78_;
  assign new_nj8_ = new_n_n822_ | new_n_n823_;
  assign new_n_n816_ = new_no0_ & new_n_n110_ & new_n_n147_;
  assign new_nv8_ = new_n_n798_ | new_n_n799_;
  assign new_n_n792_ = new_no0_ & new_n_n134_ & new_n_n147_;
  assign new_n_n785_ = new_n_n194_ & new_n_n141_ & new_n_n145_;
  assign new_ng9_ = new_n_n776_ | new_n_n777_;
  assign new_n_n761_ = new_ni4_ & new_nl4_ & new_n_n184_;
  assign new_ng15_ = new_n_n195_ | new_n_n755_ | new_n_n754_;
  assign new_nw15_ = new_n_n750_ | new_n_n748_ | new_n_n751_;
  assign new_n_n748_ = new_n_n204_ & new_n_n201_;
  assign new_nh16_ = new_n_n746_ | new_nk1_;
  assign new_n_n744_ = new_n_n208_ & new_n_n378_ & new_n_n254_;
  assign new_ni17_ = new_n_n739_ | new_n_n212_;
  assign new_n_n735_ = new_n_n217_ & new_n_n378_ & new_n_n254_;
  assign new_nu18_ = new_n_n231_ & new_nl4_;
  assign new_ng19_ = new_n_n719_ | new_n_n232_;
  assign new_n_n715_ = new_n_n237_ & new_n_n378_ & new_n_n254_;
  assign new_nb20_ = new_n_n710_ | new_n_n742_ | new_n_n697_;
  assign new_na21_ = new_n_n700_ | new_n_n742_ | new_n_n697_;
  assign new_ni21_ = new_n_n694_ | new_n_n693_ | new_n_n692_;
  assign new_n_n686_ = new_n_n428_ & new_n_n350_ & new_n_n263_;
  assign new_nf22_ = new_n_n679_ | new_n_n678_ | new_n_n677_;
  assign new_n_n677_ = new_nk0_ & new_n_n430_ & new_nl_;
  assign new_no22_ = new_no2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n666_ = new_n_n428_ & new_n_n350_ & new_n_n275_;
  assign new_nh23_ = new_n_n659_ | new_n_n658_ | new_n_n657_;
  assign new_n_n628_ = new_nl_ & new_n_n305_ & new_n_n353_;
  assign new_no24_ = new_n_n617_ | new_n_n619_ | new_n_n618_ | new_n_n620_;
  assign new_n_n618_ = new_n_n298_ & new_n_n300_ & new_n_n299_;
  assign new_nt24_ = new_nz2_ & new_nl4_;
  assign new_nb25_ = new_n_n439_ | new_n_n417_ | new_nj25_;
  assign new_ng25_ = new_nl1_ | new_nk1_ | new_nj1_;
  assign new_nm27_ = new_n_n439_ | new_n_n420_ | new_nj25_;
  assign new_nc28_ = new_nq0_ | new_n_n324_;
  assign new_nh28_ = new_n_n411_ | new_nq0_;
  assign new_n_n585_ = new_nh6_ & new_ni6_ & new_n_n329_;
  assign new_nr28_ = new_nh1_ & new_ni6_;
  assign new_n_n570_ = new_nj6_ & new_n_n337_ & new_n_n336_;
  assign new_nd30_ = new_no0_ & new_n_n432_ & new_nm0_;
  assign new_no30_ = new_n_n437_ | new_n_n458_ | new_nx3_;
  assign new_n_n543_ = new_n_n404_ & new_nl25_ & new_n_n370_;
  assign new_no31_ = new_nj25_ | new_n_n412_ | new_nq0_;
  assign new_nv31_ = new_ne4_ & new_n_n454_ & new_no4_;
  assign new_n_n519_ = new_n_n413_ & new_nl0_;
  assign new_nm33_ = new_n_n428_ & new_n_n416_;
  assign new_n_n496_ = new_n_n431_ & new_n_n430_ & new_n_n423_;
  assign new_n_n489_ = new_nk0_ & new_nl0_ & new_n_n427_;
  assign new_n_n465_ = new_nz0_ & new_na1_ & new_n_n447_;
  assign new_np35_ = new_nj1_ | new_ni1_ | new_nh1_;
  assign new_n_n432_ = ~new_nn0_;
  assign new_n_n413_ = ~new_nd3_;
  assign new_n_n382_ = ~new_ne32_;
  assign new_n_n371_ = ~new_nm31_;
  assign new_n_n316_ = ~new_nx34_;
  assign new_n_n305_ = ~new_nr23_;
  assign new_n_n283_ = ~new_no23_;
  assign new_n_n272_ = ~new_nt22_;
  assign new_n_n217_ = ~new_nr1_;
  assign new_n_n206_ = ~new_ng15_;
  assign new_n_n195_ = ~new_nh35_;
  assign new_n_n184_ = ~new_ni32_;
  assign new_n_n173_ = ~new_nh31_;
  assign new_n_n118_ = ~new_np26_;
  assign new_n_n107_ = ~new_nz25_;
  assign new_n_n96_ = ~new_nk24_;
  assign new_n_n85_ = ~new_nq21_;
  assign new_n_n9_ = ~new_ns33_;
  assign new_n_n1080_ = new_n_n431_ & new_n_n430_ & new_n_n14_;
  assign new_na5_ = new_n_n1073_ | new_n_n1072_ | new_n_n1071_;
  assign new_n_n1010_ = new_n_n41_ & new_n_n432_ & new_n_n42_;
  assign new_n_n1002_ = new_na17_ & new_n_n432_ & new_n_n44_;
  assign new_n_n923_ = new_n_n61_ & new_nz1_ & new_n_n62_;
  assign new_n_n915_ = new_na17_ & new_na2_ & new_n_n64_;
  assign new_n_n863_ = new_n_n73_ & new_n_n83_ & new_n_n74_;
  assign new_n_n855_ = new_na17_ & new_n_n83_ & new_n_n76_;
  assign new_n_n835_ = new_n_n350_ & new_n_n83_ & new_n_n80_;
  assign new_n_n823_ = new_n_n194_ & new_n_n103_ & new_n_n145_;
  assign new_n_n817_ = new_n_n194_ & new_n_n109_ & new_n_n145_;
  assign new_n_n799_ = new_n_n194_ & new_n_n127_ & new_n_n145_;
  assign new_n_n793_ = new_n_n194_ & new_n_n133_ & new_n_n145_;
  assign new_n_n784_ = new_no0_ & new_n_n142_ & new_n_n147_;
  assign new_n_n778_ = new_no0_ & new_n_n152_ & new_n_n151_;
  assign new_n_n760_ = new_nn1_ & new_nl4_ & new_n_n184_;
  assign new_nw9_ = new_n_n194_ & new_nk4_;
  assign new_n_n751_ = new_n_n204_ & new_nd1_;
  assign new_nf16_ = new_n_n750_ | new_n_n748_ | new_n_n747_;
  assign new_nj16_ = new_nc1_ | new_nn0_ | new_n_n203_;
  assign new_nv16_ = new_n_n744_ | new_n_n207_;
  assign new_n_n739_ = new_n_n213_ & new_n_n378_ & new_n_n254_;
  assign new_ns17_ = new_n_n735_ | new_n_n216_;
  assign new_nw18_ = new_n_n723_ | new_n_n228_;
  assign new_ne19_ = new_n_n235_ & new_nl4_;
  assign new_nr19_ = new_n_n714_ | new_n_n742_ | new_n_n697_;
  assign new_n_n711_ = new_n_n241_ & new_n_n378_ & new_n_n254_;
  assign new_n_n700_ = new_nb0_ & new_no0_ & new_n_n408_;
  assign new_n_n695_ = new_n_n387_ & new_n_n258_ & new_n_n279_;
  assign new_n_n685_ = new_n_n387_ & new_n_n264_ & new_n_n279_;
  assign new_n_n680_ = new_n_n387_ & new_n_n267_ & new_n_n279_;
  assign new_ng22_ = new_no2_ | new_n_n365_;
  assign new_nn22_ = new_np2_ | new_n_n365_;
  assign new_n_n665_ = new_n_n387_ & new_n_n276_ & new_n_n279_;
  assign new_n_n660_ = new_n_n387_ & new_n_n280_ & new_n_n279_;
  assign new_n_n627_ = new_n_n365_ & new_nv2_ & new_n_n306_;
  assign new_n_n621_ = new_n_n365_ & new_nw2_ & new_n_n306_;
  assign new_n_n617_ = new_n_n387_ & new_n_n300_ & new_n_n299_;
  assign new_n_n611_ = new_n_n387_ & new_n_n304_ & new_n_n303_;
  assign new_nc25_ = new_n_n309_ | new_n_n607_ | new_n_n606_;
  assign new_nf25_ = new_nj1_ | new_ni1_ | new_n_n338_;
  assign new_nn27_ = new_nq0_ | new_n_n323_;
  assign new_nb28_ = new_n_n439_ | new_n_n325_ | new_nj25_;
  assign new_ni28_ = new_n_n439_ | new_nj25_ | new_n_n412_;
  assign new_nl28_ = new_n_n582_ | new_n_n584_ | new_n_n583_ | new_n_n585_;
  assign new_ns28_ = new_n_n577_ | new_n_n578_;
  assign new_n_n571_ = new_n_n400_ & new_n_n337_ & new_n_n336_;
  assign new_ne30_ = new_nx3_ | new_n_n458_;
  assign new_nn30_ = new_no0_ & new_n_n432_ & new_n_n428_;
  assign new_nt30_ = new_nq0_ | new_ng1_;
  assign new_np31_ = new_n_n456_ | new_ng1_ | new_nq0_;
  assign new_nu31_ = new_n_n439_ | new_n_n460_ | new_n_n461_;
  assign new_n_n518_ = new_n_n429_ & new_n_n430_;
  assign new_n_n512_ = new_n_n427_ & new_n_n415_;
  assign new_nw33_ = new_n_n428_ | new_n_n495_ | new_n_n494_;
  assign new_nz33_ = new_n_n428_ | new_n_n489_ | new_n_n488_;
  assign new_ni35_ = new_n_n460_ | new_n_n461_ | new_n_n448_;
  assign new_no35_ = new_ng4_ | new_nh4_;
  assign new_nl6_ = ~new_nl1_;
  assign new_n_n403_ = ~new_nx32_;
  assign new_n_n381_ = ~new_nd32_;
  assign new_n_n372_ = ~new_nj31_;
  assign new_n_n315_ = ~new_nm25_;
  assign new_n_n306_ = ~new_nt23_;
  assign new_n_n282_ = ~new_nq23_;
  assign new_n_n273_ = ~new_nu22_;
  assign new_n_n216_ = ~new_nt17_;
  assign new_n_n207_ = ~new_nx16_;
  assign new_n_n185_ = ~new_nj28_;
  assign new_n_n183_ = ~new_nz31_;
  assign new_n_n174_ = ~new_nr31_;
  assign new_n_n117_ = ~new_no26_;
  assign new_n_n108_ = ~new_na26_;
  assign new_n_n95_ = ~new_ng24_;
  assign new_n_n86_ = ~new_nx21_;
  assign new_nx4_ = new_n_n1082_ | new_n_n1081_ | new_n_n1080_;
  assign new_n_n1074_ = new_n_n431_ & new_n_n430_ & new_n_n16_;
  assign new_n_n1013_ = new_n_n41_ & new_np1_ & new_n_n42_;
  assign new_n_n1003_ = new_n_n350_ & new_nq1_ & new_n_n44_;
  assign new_nj7_ = new_n_n914_ | new_n_n912_ | new_n_n911_ | new_n_n913_ | new_n_n915_ | new_n_n910_ | new_n_n909_ | new_n_n908_ | new_n_n907_;
  assign new_n_n862_ = new_n_n350_ & new_n_n83_ & new_n_n74_;
  assign new_n_n846_ = new_na17_ & new_n_n83_ & new_n_n78_;
  assign new_n_n836_ = new_n_n79_ & new_n_n83_ & new_n_n80_;
  assign new_n_n810_ = new_no0_ & new_n_n116_ & new_n_n147_;
  assign new_n_n803_ = new_n_n194_ & new_n_n123_ & new_n_n145_;
  assign new_n_n798_ = new_no0_ & new_n_n128_ & new_n_n147_;
  assign new_n_n791_ = new_n_n194_ & new_n_n135_ & new_n_n145_;
  assign new_n_n786_ = new_no0_ & new_n_n140_ & new_n_n147_;
  assign new_n_n779_ = new_n_n150_ & new_n_n149_ & new_n_n185_;
  assign new_ns9_ = new_n_n758_ | new_n_n759_;
  assign new_n_n754_ = new_n_n317_ & new_ni1_ & new_n_n196_;
  assign new_n_n752_ = new_nc1_ & new_ne1_;
  assign new_nd16_ = new_n_n746_ | new_nj1_;
  assign new_nl16_ = new_nq0_ | new_n_n411_ | new_n_n746_;
  assign new_n_n743_ = new_nj0_ & new_no0_ & new_n_n408_;
  assign new_n_n740_ = new_ni0_ & new_no0_ & new_n_n408_;
  assign new_nq17_ = new_n_n219_ & new_nl4_;
  assign new_n_n723_ = new_n_n229_ & new_n_n378_ & new_n_n254_;
  assign new_nh19_ = new_n_n718_ | new_n_n742_ | new_n_n697_;
  assign new_no19_ = new_n_n239_ & new_nl4_;
  assign new_na20_ = new_n_n711_ | new_n_n240_;
  assign new_ng20_ = new_n_n708_ | new_n_n742_ | new_n_n697_;
  assign new_n_n704_ = new_nz_ & new_no0_ & new_n_n408_;
  assign new_nt21_ = new_nl2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n681_ = new_n_n428_ & new_n_n350_ & new_n_n266_;
  assign new_nh22_ = new_nn2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n671_ = new_n_n428_ & new_n_n350_ & new_n_n272_;
  assign new_nv22_ = new_np2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n661_ = new_n_n428_ & new_n_n350_ & new_n_n278_;
  assign new_nh24_ = new_nw2_ & new_nl4_;
  assign new_n_n622_ = new_nm_ & new_n_n305_ & new_n_n353_;
  assign new_np24_ = new_ny2_ & new_nl4_;
  assign new_n_n610_ = new_no_ & new_n_n305_ & new_n_n353_;
  assign new_n_n608_ = new_n_n428_ & new_n_n350_ & new_n_n353_;
  assign new_n_n602_ = new_n_n330_ & new_n_n335_ & new_n_n311_;
  assign new_nj27_ = new_n_n439_ | new_n_n323_ | new_nj25_;
  assign new_nz27_ = new_nq0_ | new_n_n414_;
  assign new_nj28_ = new_n_n590_ | new_n_n588_ | new_n_n587_ | new_n_n586_ | new_n_n589_ | new_n_n591_;
  assign new_n_n583_ = new_nh6_ & new_n_n335_ & new_n_n329_;
  assign new_n_n579_ = new_ni6_ & new_nh6_ & new_n_n335_;
  assign new_n_n572_ = new_nj1_ & new_n_n338_ & new_n_n336_;
  assign new_n_n547_ = new_n_n387_ & new_n_n359_ & new_n_n358_;
  assign new_nm30_ = new_n_n378_ | new_nq0_ | new_n_n364_;
  assign new_nu30_ = new_n_n544_ | new_n_n545_;
  assign new_nf31_ = new_nd4_ | new_n_n439_;
  assign new_n_n539_ = new_nk0_ & new_n_n430_ & new_nm0_;
  assign new_n_n520_ = new_n_n429_ & new_nl0_;
  assign new_n_n513_ = new_n_n427_ & new_n_n430_;
  assign new_n_n509_ = new_n_n417_ & new_nl0_;
  assign new_ns33_ = new_n_n428_ & new_n_n420_;
  assign new_n_n467_ = new_nk6_ & new_nz0_ & new_n_n447_;
  assign new_nn35_ = new_n_n456_ & new_n_n457_;
  assign new_n_n448_ = ~new_nn35_;
  assign new_n_n394_ = ~new_nv0_;
  assign new_n_n384_ = ~new_nc32_;
  assign new_n_n373_ = ~new_nl31_;
  assign new_n_n296_ = ~new_nm24_;
  assign new_n_n285_ = ~new_nu23_;
  assign new_n_n274_ = ~new_nc23_;
  assign new_n_n215_ = ~new_nq1_;
  assign new_n_n197_ = ~new_no15_;
  assign new_n_n186_ = ~new_nl32_;
  assign new_n_n116_ = ~new_nm26_;
  assign new_n_n105_ = ~new_nw25_;
  assign new_n_n98_ = ~new_ns24_;
  assign new_n_n87_ = ~new_ne22_;
  assign new_n_n1082_ = new_n_n14_ & new_no3_;
  assign new_n_n1075_ = new_nk0_ & new_nl0_ & new_n_n16_;
  assign new_n_n1012_ = new_n_n350_ & new_np1_ & new_n_n42_;
  assign new_n_n1004_ = new_n_n43_ & new_nq1_ & new_n_n44_;
  assign new_ni7_ = new_n_n923_ | new_n_n921_ | new_n_n920_ | new_n_n922_ | new_n_n924_ | new_n_n919_ | new_n_n918_ | new_n_n917_ | new_n_n916_;
  assign new_n_n853_ = new_n_n350_ & new_n_n83_ & new_n_n76_;
  assign new_n_n845_ = new_n_n77_ & new_n_n83_ & new_n_n78_;
  assign new_n_n837_ = new_na17_ & new_n_n83_ & new_n_n80_;
  assign new_nq8_ = new_n_n808_ | new_n_n809_;
  assign new_nt8_ = new_n_n802_ | new_n_n803_;
  assign new_nw8_ = new_n_n796_ | new_n_n797_;
  assign new_nz8_ = new_n_n790_ | new_n_n791_;
  assign new_nc9_ = new_n_n784_ | new_n_n785_;
  assign new_nf9_ = new_n_n778_ | new_n_n779_;
  assign new_n_n759_ = new_n_n187_ & new_n_n186_ & new_n_n185_;
  assign new_n_n755_ = new_n_n410_ & new_nh1_ & new_n_n196_;
  assign new_nt15_ = new_nl6_ & new_nk6_ & new_n_n198_;
  assign new_nc16_ = new_nq0_ | new_n_n411_ | new_n_n200_;
  assign new_n_n746_ = new_n_n432_ & new_n_n204_ & new_nt15_;
  assign new_nx16_ = new_n_n743_ | new_n_n742_ | new_n_n697_;
  assign new_ng17_ = new_n_n215_ & new_nl4_;
  assign new_n_n736_ = new_ng0_ & new_no0_ & new_n_n408_;
  assign new_nx18_ = new_n_n722_ | new_n_n742_ | new_n_n697_;
  assign new_n_n719_ = new_n_n233_ & new_n_n378_ & new_n_n254_;
  assign new_nq19_ = new_n_n715_ | new_n_n236_;
  assign new_ny19_ = new_n_n243_ & new_nl4_;
  assign new_n_n708_ = new_nx_ & new_no0_ & new_n_n408_;
  assign new_nq20_ = new_n_n704_ | new_n_n742_ | new_n_n697_;
  assign new_nx21_ = new_n_n262_ | new_n_n686_ | new_n_n685_;
  assign new_ne22_ = new_n_n265_ | new_n_n681_ | new_n_n680_;
  assign new_nl22_ = new_n_n268_ | new_n_n676_ | new_n_n675_;
  assign new_ns22_ = new_n_n271_ | new_n_n671_ | new_n_n670_;
  assign new_nz22_ = new_n_n274_ | new_n_n666_ | new_n_n665_;
  assign new_ng23_ = new_n_n277_ | new_n_n661_ | new_n_n660_;
  assign new_ni24_ = new_n_n627_ | new_n_n628_;
  assign new_nm24_ = new_n_n621_ | new_n_n622_;
  assign new_nq24_ = new_n_n615_ | new_n_n616_;
  assign new_nu24_ = new_n_n609_ | new_n_n610_;
  assign new_na25_ = new_n_n412_ | new_nq0_ | new_n_n411_;
  assign new_n_n603_ = new_nh6_ & new_n_n335_ & new_n_n311_;
  assign new_nk27_ = new_nq0_ | new_n_n322_;
  assign new_ny27_ = new_n_n439_ | new_n_n324_ | new_nj25_;
  assign new_n_n591_ = new_nh1_ & new_n_n395_;
  assign new_n_n584_ = new_n_n330_ & new_ni6_ & new_n_n329_;
  assign new_nq28_ = new_n_n529_ | new_nj6_;
  assign new_n_n573_ = new_n_n393_ & new_n_n338_ & new_n_n336_;
  assign new_nc30_ = new_n_n378_ | new_nq0_ | new_n_n360_;
  assign new_n_n546_ = new_n_n387_ & new_n_n363_ & new_n_n362_;
  assign new_n_n545_ = new_n_n366_ & new_n_n454_;
  assign new_ne31_ = new_n_n439_ | new_ne4_ | new_nd4_;
  assign new_nn31_ = new_n_n411_ | new_n_n374_ | new_n_n375_;
  assign new_ni33_ = new_n_n519_ | new_n_n518_ | new_n_n517_;
  assign new_n_n514_ = new_n_n415_ & new_nl0_;
  assign new_n_n508_ = new_n_n426_ & new_n_n430_;
  assign new_n_n502_ = new_n_n425_ & new_n_n419_;
  assign new_n_n466_ = new_nj6_ & new_na1_ & new_n_n447_;
  assign new_nm35_ = new_ne4_ & new_nf4_;
  assign new_n_n458_ = ~new_ny3_;
  assign new_n_n385_ = ~new_nb32_;
  assign new_n_n383_ = ~new_nf32_;
  assign new_n_n374_ = ~new_nv31_;
  assign new_n_n295_ = ~new_nw2_;
  assign new_n_n286_ = ~new_nt2_;
  assign new_n_n284_ = ~new_nw23_;
  assign new_n_n205_ = ~new_nd1_;
  assign new_n_n196_ = ~new_ng35_;
  assign new_n_n187_ = ~new_nk32_;
  assign new_n_n115_ = ~new_nl26_;
  assign new_n_n106_ = ~new_nx25_;
  assign new_n_n97_ = ~new_no24_;
  assign new_n_n88_ = ~new_nl22_;
  assign new_nc5_ = new_n_n1067_ | new_n_n1066_ | new_n_n1065_;
  assign new_nk5_ = new_nm0_ & new_nt3_;
  assign new_n_n1057_ = new_n_n436_ & new_n_n435_;
  assign new_n_n1050_ = new_nn0_ & new_n_n32_ & new_n_n27_;
  assign new_n_n1041_ = new_nn0_ & new_no4_ & new_n_n31_;
  assign new_n_n995_ = new_n_n45_ & new_nr1_ & new_n_n46_;
  assign new_n_n985_ = new_n_n350_ & new_ns1_ & new_n_n48_;
  assign new_n_n975_ = new_na17_ & new_n_n432_ & new_n_n50_;
  assign new_n_n965_ = new_n_n51_ & new_n_n432_ & new_n_n52_;
  assign new_n_n955_ = new_n_n350_ & new_n_n432_ & new_n_n54_;
  assign new_n_n945_ = new_na17_ & new_n_n83_ & new_n_n56_;
  assign new_n_n935_ = new_n_n57_ & new_n_n83_ & new_n_n58_;
  assign new_n_n925_ = new_n_n350_ & new_n_n83_ & new_n_n60_;
  assign new_nl7_ = new_n_n896_ | new_n_n894_ | new_n_n893_ | new_n_n895_ | new_n_n897_ | new_n_n892_ | new_n_n891_ | new_n_n890_ | new_n_n889_;
  assign new_n_n888_ = new_na17_ & new_nd2_ & new_n_n70_;
  assign new_n_n878_ = new_n_n71_ & new_ne2_ & new_n_n72_;
  assign new_n_n868_ = new_n_n350_ & new_nf2_ & new_n_n74_;
  assign new_n_n858_ = new_na17_ & new_n_n432_ & new_n_n76_;
  assign new_n_n848_ = new_n_n77_ & new_n_n432_ & new_n_n78_;
  assign new_n_n838_ = new_n_n350_ & new_n_n432_ & new_n_n80_;
  assign new_n_n802_ = new_no0_ & new_n_n124_ & new_n_n147_;
  assign new_n_n795_ = new_n_n194_ & new_n_n131_ & new_n_n145_;
  assign new_nb9_ = new_n_n786_ | new_n_n787_;
  assign new_n_n780_ = new_no0_ & new_n_n148_ & new_n_n147_;
  assign new_n_n772_ = new_no0_ & new_n_n161_ & new_n_n160_;
  assign new_np9_ = new_n_n174_ | new_n_n765_ | new_n_n764_;
  assign new_no17_ = new_n_n736_ | new_n_n742_ | new_n_n697_;
  assign new_n_n731_ = new_n_n221_ & new_n_n378_ & new_n_n254_;
  assign new_nn18_ = new_n_n726_ | new_n_n742_ | new_n_n697_;
  assign new_n_n655_ = new_n_n428_ & new_n_n432_ & new_nt15_;
  assign new_nr23_ = new_n_n378_ | new_nn0_ | new_nm0_;
  assign new_n_n643_ = new_n_n286_ & new_na17_ & new_n_n287_;
  assign new_n_n635_ = new_n_n387_ & new_n_n291_ & new_n_n290_;
  assign new_n_n599_ = new_nj1_ & new_nk1_;
  assign new_n_n595_ = new_n_n319_ & new_n_n396_;
  assign new_nd26_ = new_nq0_ | new_n_n413_;
  assign new_nu26_ = new_n_n439_ | new_n_n427_ | new_nj25_;
  assign new_nb29_ = new_n_n697_ | new_n_n742_;
  assign new_nk29_ = new_nl4_ & new_n_n437_ & new_n_n345_;
  assign new_n_n556_ = new_n_n347_ & new_n_n349_ & new_n_n348_;
  assign new_nt29_ = new_n_n548_ | new_n_n549_;
  assign new_nh30_ = new_nl4_ & new_n_n433_ & new_n_n441_;
  assign new_n_n536_ = new_nh6_ & new_n_n389_ & new_n_n390_;
  assign new_nr32_ = new_n_n397_ | new_n_n528_ | new_n_n527_;
  assign new_ny32_ = new_nn4_ & new_nk4_ & new_n_n405_;
  assign new_nk33_ = new_n_n516_ | new_n_n515_ | new_n_n512_;
  assign new_no33_ = new_n_n509_ | new_n_n508_ | new_n_n507_;
  assign new_n_n482_ = new_nj6_ & new_na1_ & new_nb1_;
  assign new_n_n472_ = new_ny0_ & new_nz0_ & new_n_n442_;
  assign new_n_n463_ = new_n_n451_ & new_n_n450_;
  assign new_n_n460_ = ~new_nf4_;
  assign new_n_n449_ = ~new_nn4_;
  assign new_n_n393_ = ~new_nw0_;
  assign new_n_n378_ = ~new_nt15_;
  assign new_n_n367_ = ~new_nw30_;
  assign new_n_n356_ = ~new_ng30_;
  assign new_n_n345_ = ~new_nl29_;
  assign new_n_n279_ = ~new_nk21_;
  assign new_n_n268_ = ~new_no22_;
  assign new_n_n257_ = ~new_ni21_;
  assign new_n_n246_ = ~new_nq20_;
  assign new_n_n235_ = ~new_na2_;
  assign new_n_n180_ = ~new_nz29_;
  assign new_n_n169_ = ~new_nv30_;
  assign new_n_n158_ = ~new_nn29_;
  assign new_n_n147_ = ~new_ne25_;
  assign new_n_n136_ = ~new_nq27_;
  assign new_n_n125_ = ~new_na27_;
  assign new_n_n5_ = ~new_nk33_;
  assign new_n_n1067_ = new_n_n19_ & new_nt3_;
  assign new_nj5_ = new_nm0_ & new_ns3_;
  assign new_no6_ = new_n_n434_ & new_n_n433_ & new_n_n22_;
  assign new_n_n1051_ = new_n_n378_ & new_n_n32_ & new_n_n27_;
  assign new_n_n1033_ = new_n_n432_ & new_np0_ & new_n_n36_;
  assign new_n_n994_ = new_n_n350_ & new_nr1_ & new_n_n46_;
  assign new_n_n986_ = new_n_n47_ & new_ns1_ & new_n_n48_;
  assign new_n_n974_ = new_n_n49_ & new_n_n432_ & new_n_n50_;
  assign new_n_n966_ = new_na17_ & new_n_n432_ & new_n_n52_;
  assign new_n_n954_ = new_na17_ & new_n_n83_ & new_n_n54_;
  assign new_n_n946_ = new_n_n350_ & new_n_n432_ & new_n_n56_;
  assign new_n_n934_ = new_n_n350_ & new_n_n83_ & new_n_n58_;
  assign new_n_n926_ = new_n_n59_ & new_n_n83_ & new_n_n60_;
  assign new_nk7_ = new_n_n905_ | new_n_n903_ | new_n_n902_ | new_n_n904_ | new_n_n906_ | new_n_n901_ | new_n_n900_ | new_n_n899_ | new_n_n898_;
  assign new_n_n887_ = new_n_n69_ & new_nd2_ & new_n_n70_;
  assign new_n_n879_ = new_na17_ & new_ne2_ & new_n_n72_;
  assign new_n_n867_ = new_na17_ & new_n_n432_ & new_n_n74_;
  assign new_n_n859_ = new_n_n350_ & new_ng2_ & new_n_n76_;
  assign new_n_n847_ = new_n_n350_ & new_n_n432_ & new_n_n78_;
  assign new_n_n839_ = new_n_n79_ & new_n_n432_ & new_n_n80_;
  assign new_nu8_ = new_n_n800_ | new_n_n801_;
  assign new_nx8_ = new_n_n794_ | new_n_n795_;
  assign new_n_n787_ = new_n_n194_ & new_n_n139_ & new_n_n145_;
  assign new_n_n781_ = new_n_n194_ & new_n_n146_ & new_n_n145_;
  assign new_nl9_ = new_n_n162_ | new_n_n771_ | new_n_n770_;
  assign new_n_n766_ = new_n_n173_ & new_nf4_;
  assign new_ne17_ = new_n_n740_ | new_n_n742_ | new_n_n697_;
  assign new_nd18_ = new_n_n730_ | new_n_n742_ | new_n_n697_;
  assign new_n_n727_ = new_n_n225_ & new_n_n378_ & new_n_n254_;
  assign new_nn23_ = new_n_n651_ | new_n_n653_ | new_n_n652_ | new_n_n654_;
  assign new_n_n649_ = new_n_n365_ & new_ns2_ & new_n_n306_;
  assign new_n_n642_ = new_n_n286_ & new_n_n288_ & new_n_n287_;
  assign new_n_n636_ = new_n_n289_ & new_n_n291_ & new_n_n290_;
  assign new_nl25_ = new_n_n316_ | new_n_n523_ | new_n_n598_;
  assign new_n_n596_ = new_n_n319_ & new_nh1_;
  assign new_nf26_ = new_n_n439_ | new_n_n422_ | new_nj25_;
  assign new_ns26_ = new_nq0_ | new_n_n425_;
  assign new_nd29_ = new_nl4_ & new_n_n440_ & new_n_n387_;
  assign new_n_n564_ = new_nn0_ & new_n_n408_ & new_n_n344_;
  assign new_n_n555_ = new_n_n350_ & new_n_n349_ & new_n_n348_;
  assign new_n_n550_ = new_nt15_ & new_n_n353_ & new_n_n352_;
  assign new_nr30_ = new_nl4_ & new_n_n434_ & new_n_n433_;
  assign new_nd32_ = new_n_n404_ & new_no4_;
  assign new_n_n528_ = new_n_n398_ & new_ni1_;
  assign new_n_n524_ = new_nk6_ & new_nl6_ & new_n_n404_;
  assign new_n_n516_ = new_n_n415_ & new_n_n430_;
  assign new_n_n510_ = new_n_n426_ & new_nl0_;
  assign new_n_n481_ = new_nz0_ & new_nk6_ & new_nb1_;
  assign new_n_n473_ = new_ni6_ & new_nz0_ & new_n_n442_;
  assign new_n_n462_ = new_n_n452_ & new_nl1_ & new_n_n451_;
  assign new_n_n461_ = ~new_ne4_;
  assign new_ni6_ = ~new_ni1_;
  assign new_n_n402_ = ~new_nw32_;
  assign new_n_n377_ = ~new_nk31_;
  assign new_n_n368_ = ~new_nf31_;
  assign new_n_n355_ = ~new_nu29_;
  assign new_n_n346_ = ~new_no29_;
  assign new_n_n278_ = ~new_nh23_;
  assign new_n_n269_ = ~new_nm22_;
  assign new_n_n256_ = ~new_nl21_;
  assign new_n_n247_ = ~new_ng2_;
  assign new_n_n225_ = ~new_nv1_;
  assign new_n_n179_ = ~new_nc30_;
  assign new_n_n170_ = ~new_nc31_;
  assign new_n_n157_ = ~new_ni29_;
  assign new_n_n148_ = ~new_nf28_;
  assign new_n_n135_ = ~new_np27_;
  assign new_n_n126_ = ~new_nb27_;
  assign new_n_n6_ = ~new_np33_;
  assign new_n_n1066_ = new_nk0_ & new_nl0_ & new_n_n19_;
  assign new_nw5_ = new_n_n1063_ | new_n_n1061_ | new_n_n1060_ | new_n_n1059_ | new_n_n1062_ | new_n_n1064_;
  assign new_nn6_ = new_n_n1057_ | new_n_n1058_;
  assign new_n_n1052_ = new_n_n28_ & new_no4_ & new_n_n27_;
  assign new_n_n1024_ = new_n_n350_ & new_n_n83_ & new_n_n38_;
  assign new_n_n993_ = new_na17_ & new_n_n432_ & new_n_n46_;
  assign new_n_n983_ = new_n_n47_ & new_n_n432_ & new_n_n48_;
  assign new_n_n977_ = new_n_n49_ & new_nt1_ & new_n_n50_;
  assign new_n_n967_ = new_n_n350_ & new_nu1_ & new_n_n52_;
  assign new_n_n953_ = new_n_n53_ & new_n_n83_ & new_n_n54_;
  assign new_n_n943_ = new_n_n350_ & new_n_n83_ & new_n_n56_;
  assign new_n_n937_ = new_n_n350_ & new_n_n432_ & new_n_n58_;
  assign new_n_n927_ = new_na17_ & new_n_n83_ & new_n_n60_;
  assign new_n_n906_ = new_na17_ & new_nb2_ & new_n_n66_;
  assign new_n_n896_ = new_n_n67_ & new_nc2_ & new_n_n68_;
  assign new_nn7_ = new_n_n878_ | new_n_n876_ | new_n_n875_ | new_n_n877_ | new_n_n879_ | new_n_n874_ | new_n_n873_ | new_n_n872_ | new_n_n871_;
  assign new_n_n866_ = new_n_n73_ & new_n_n432_ & new_n_n74_;
  assign new_n_n856_ = new_n_n350_ & new_n_n432_ & new_n_n76_;
  assign new_n_n850_ = new_n_n350_ & new_nh2_ & new_n_n78_;
  assign new_n_n840_ = new_na17_ & new_n_n432_ & new_n_n80_;
  assign new_n_n827_ = new_n_n81_ & new_n_n83_ & new_n_n82_;
  assign new_nc8_ = new_n_n408_ & new_no0_ & new_n_n93_;
  assign new_n_n801_ = new_n_n194_ & new_n_n125_ & new_n_n145_;
  assign new_ny8_ = new_n_n792_ | new_n_n793_;
  assign new_n_n789_ = new_n_n194_ & new_n_n137_ & new_n_n145_;
  assign new_ne9_ = new_n_n780_ | new_n_n781_;
  assign new_nk9_ = new_n_n179_ | new_n_n773_ | new_n_n772_;
  assign new_no9_ = new_n_n411_ | new_n_n172_ | new_n_n766_;
  assign new_nu16_ = new_na17_ | new_n_n365_;
  assign new_na18_ = new_n_n223_ & new_nl4_;
  assign new_nm18_ = new_n_n727_ | new_n_n224_;
  assign new_n_n654_ = new_n_n282_ & new_n_n301_;
  assign new_nt23_ = new_n_n432_ & new_n_n428_ & new_n_n285_;
  assign new_ny23_ = new_n_n641_ | new_n_n643_ | new_n_n642_ | new_n_n644_;
  assign new_n_n637_ = new_n_n289_ & new_na17_ & new_n_n290_;
  assign new_nk24_ = new_n_n623_ | new_n_n625_ | new_n_n624_ | new_n_n626_;
  assign new_n_n598_ = new_n_n317_ & new_ni1_;
  assign new_n_n594_ = new_nk1_ & new_nj1_;
  assign new_na26_ = new_nq0_ | new_n_n415_;
  assign new_nr26_ = new_n_n439_ | new_n_n426_ | new_nj25_;
  assign new_np27_ = new_n_n439_ | new_n_n418_ | new_nj25_;
  assign new_nf28_ = new_nq0_ | new_n_n325_;
  assign new_ne29_ = new_n_n566_ | new_n_n567_;
  assign new_nm29_ = new_n_n458_ | new_n_n365_;
  assign new_n_n558_ = new_n_n350_ & new_n_n432_ & new_n_n348_;
  assign new_n_n551_ = new_na4_ & new_n_n353_ & new_n_n352_;
  assign new_nf30_ = new_n_n365_ | new_na4_ | new_n_n437_;
  assign new_nq30_ = new_n_n441_ & new_nz3_ & new_ny3_;
  assign new_ne32_ = new_nf4_ & new_ne4_ & new_n_n454_;
  assign new_n_n534_ = new_nh1_ & new_n_n391_ & new_n_n390_;
  assign new_n_n525_ = new_n_n404_ & new_nj6_;
  assign new_n_n517_ = new_n_n429_ & new_n_n413_;
  assign new_n_n511_ = new_n_n417_ & new_n_n430_;
  assign new_nf34_ = new_n_n439_ & new_nl1_ & new_n_n432_;
  assign new_np34_ = new_nh1_ & new_nl4_;
  assign new_nj35_ = new_n_n464_ | new_n_n463_ | new_n_n462_;
  assign new_nr35_ = new_ng4_ | new_n_n460_ | new_n_n461_;
  assign new_n_n433_ = ~new_nb4_;
  assign new_n_n412_ = ~new_nl25_;
  assign new_n_n380_ = ~new_nt31_;
  assign new_n_n369_ = ~new_nd31_;
  assign new_n_n336_ = ~new_nw28_;
  assign new_n_n325_ = ~new_nv3_;
  assign new_n_n281_ = ~new_ns2_;
  assign new_n_n270_ = ~new_nn22_;
  assign new_n_n255_ = ~new_nj2_;
  assign new_n_n237_ = ~new_nb2_;
  assign new_n_n226_ = ~new_ns18_;
  assign new_n_n182_ = ~new_na32_;
  assign new_n_n171_ = ~new_nb31_;
  assign new_n_n156_ = ~new_nj29_;
  assign new_n_n145_ = ~new_nc25_;
  assign new_n_n138_ = ~new_nt27_;
  assign new_n_n127_ = ~new_nd27_;
  assign new_n_n7_ = ~new_no33_;
  assign new_n_n1065_ = new_n_n431_ & new_n_n430_ & new_n_n19_;
  assign new_nl5_ = new_ng1_ & new_n_n405_;
  assign new_n_n1058_ = new_ni4_ & new_nf1_;
  assign new_n_n1053_ = new_nn0_ & new_no4_ & new_n_n27_;
  assign new_n_n1015_ = new_n_n350_ & new_n_n83_ & new_n_n40_;
  assign new_n_n992_ = new_n_n45_ & new_n_n432_ & new_n_n46_;
  assign new_n_n984_ = new_na17_ & new_n_n432_ & new_n_n48_;
  assign new_n_n976_ = new_n_n350_ & new_nt1_ & new_n_n50_;
  assign new_n_n968_ = new_n_n51_ & new_nu1_ & new_n_n52_;
  assign new_n_n952_ = new_n_n350_ & new_n_n83_ & new_n_n54_;
  assign new_n_n944_ = new_n_n55_ & new_n_n83_ & new_n_n56_;
  assign new_n_n936_ = new_na17_ & new_n_n83_ & new_n_n58_;
  assign new_n_n928_ = new_n_n350_ & new_n_n432_ & new_n_n60_;
  assign new_n_n905_ = new_n_n65_ & new_nb2_ & new_n_n66_;
  assign new_n_n897_ = new_na17_ & new_nc2_ & new_n_n68_;
  assign new_nm7_ = new_n_n887_ | new_n_n885_ | new_n_n884_ | new_n_n886_ | new_n_n888_ | new_n_n883_ | new_n_n882_ | new_n_n881_ | new_n_n880_;
  assign new_n_n865_ = new_n_n350_ & new_n_n432_ & new_n_n74_;
  assign new_n_n857_ = new_n_n75_ & new_n_n432_ & new_n_n76_;
  assign new_n_n849_ = new_na17_ & new_n_n432_ & new_n_n78_;
  assign new_n_n841_ = new_n_n350_ & new_ni2_ & new_n_n80_;
  assign new_n_n826_ = new_n_n350_ & new_n_n83_ & new_n_n82_;
  assign new_nb8_ = new_n_n408_ & new_no0_ & new_n_n92_;
  assign new_n_n800_ = new_no0_ & new_n_n126_ & new_n_n147_;
  assign new_n_n794_ = new_no0_ & new_n_n132_ & new_n_n147_;
  assign new_n_n788_ = new_no0_ & new_n_n138_ & new_n_n147_;
  assign new_n_n782_ = new_no0_ & new_n_n144_ & new_n_n147_;
  assign new_n_n773_ = new_n_n159_ & new_n_n163_ & new_n_n180_;
  assign new_n_n767_ = new_n_n171_ & new_ne4_;
  assign new_ng16_ = new_nq0_ | new_n_n411_ | new_n_n202_;
  assign new_nc18_ = new_n_n731_ | new_n_n220_;
  assign new_nk18_ = new_n_n227_ & new_nl4_;
  assign new_n_n653_ = new_n_n281_ & new_na17_ & new_n_n282_;
  assign new_ns23_ = new_n_n647_ | new_n_n648_;
  assign new_n_n644_ = new_n_n287_ & new_n_n301_;
  assign new_n_n638_ = new_n_n290_ & new_n_n301_;
  assign new_n_n620_ = new_n_n299_ & new_n_n301_;
  assign new_nm25_ = new_nl1_ | new_nk1_ | new_n_n318_;
  assign new_ns25_ = new_n_n594_ | new_n_n593_ | new_n_n592_;
  assign new_nc26_ = new_n_n439_ | new_n_n421_ | new_nj25_;
  assign new_np26_ = new_nq0_ | new_n_n424_;
  assign new_nq27_ = new_nq0_ | new_n_n420_;
  assign new_ne28_ = new_n_n439_ | new_n_n328_ | new_nj25_;
  assign new_n_n567_ = new_n_n378_ & new_n_n408_ & new_n_n341_;
  assign new_nl29_ = new_n_n458_ | new_nx3_ | new_na17_;
  assign new_n_n557_ = new_n_n346_ & new_n_n349_ & new_n_n348_;
  assign new_n_n552_ = new_na4_ & new_n_n378_ & new_n_n352_;
  assign new_ng30_ = new_ny3_ & new_nz3_;
  assign new_np30_ = new_n_n365_ | new_nb4_ | new_na4_;
  assign new_nf32_ = new_nk4_ & new_n_n457_ & new_n_n456_;
  assign new_n_n535_ = new_nh6_ & new_n_n392_ & new_n_n390_;
  assign new_nq32_ = new_ni1_ | new_n_n395_ | new_n_n396_;
  assign new_nj33_ = new_n_n428_ & new_n_n414_;
  assign new_nn33_ = new_n_n511_ | new_n_n510_ | new_n_n507_;
  assign new_ng34_ = new_n_n434_ & new_n_n433_ & new_n_n441_;
  assign new_no34_ = new_n_n439_ & new_nm1_ & new_nl1_;
  assign new_n_n464_ = new_n_n451_ & new_n_n449_;
  assign new_nq35_ = new_n_n458_ | new_nx3_ | new_n_n459_;
  assign new_n_n423_ = ~new_ng3_;
  assign new_n_n422_ = ~new_nf3_;
  assign new_n_n379_ = ~new_ns31_;
  assign new_n_n370_ = ~new_ne31_;
  assign new_n_n335_ = ~new_ng25_;
  assign new_n_n326_ = ~new_nr28_;
  assign new_n_n280_ = ~new_ni23_;
  assign new_n_n271_ = ~new_nv22_;
  assign new_n_n245_ = ~new_nf2_;
  assign new_n_n236_ = ~new_nr19_;
  assign new_n_n227_ = ~new_nw1_;
  assign new_n_n181_ = ~new_ny31_;
  assign new_n_n172_ = ~new_ni31_;
  assign new_n_n155_ = ~new_nd29_;
  assign new_n_n146_ = ~new_ne28_;
  assign new_n_n137_ = ~new_ns27_;
  assign new_n_n128_ = ~new_ne27_;
  assign new_n_n8_ = ~new_nn33_;
  assign new_n_n1103_ = new_n_n431_ & new_n_n2_ & new_n_n0_;
  assign new_nd5_ = new_nm0_ & new_nm3_;
  assign new_n_n1044_ = new_nn0_ & new_n_n32_ & new_n_n29_;
  assign new_n_n1035_ = new_no4_ & new_nl1_ & new_n_n35_;
  assign new_n_n1026_ = new_na17_ & new_n_n83_ & new_n_n38_;
  assign new_n_n1016_ = new_n_n39_ & new_n_n83_ & new_n_n40_;
  assign new_n_n991_ = new_n_n350_ & new_n_n432_ & new_n_n46_;
  assign new_n_n981_ = new_na17_ & new_n_n83_ & new_n_n48_;
  assign new_n_n971_ = new_n_n49_ & new_n_n83_ & new_n_n50_;
  assign new_n_n961_ = new_n_n350_ & new_n_n83_ & new_n_n52_;
  assign new_n_n959_ = new_n_n53_ & new_nv1_ & new_n_n54_;
  assign new_n_n949_ = new_n_n350_ & new_nw1_ & new_n_n56_;
  assign new_n_n939_ = new_na17_ & new_n_n432_ & new_n_n58_;
  assign new_n_n929_ = new_n_n59_ & new_n_n432_ & new_n_n60_;
  assign new_n_n916_ = new_n_n350_ & new_n_n83_ & new_n_n62_;
  assign new_n_n904_ = new_n_n350_ & new_nb2_ & new_n_n66_;
  assign new_n_n894_ = new_na17_ & new_n_n432_ & new_n_n68_;
  assign new_n_n884_ = new_n_n69_ & new_n_n432_ & new_n_n70_;
  assign new_n_n874_ = new_n_n350_ & new_n_n432_ & new_n_n72_;
  assign new_np7_ = new_n_n860_ | new_n_n858_ | new_n_n857_ | new_n_n859_ | new_n_n861_ | new_n_n856_ | new_n_n855_ | new_n_n854_ | new_n_n853_;
  assign new_n_n852_ = new_na17_ & new_nh2_ & new_n_n78_;
  assign new_n_n842_ = new_n_n79_ & new_ni2_ & new_n_n80_;
  assign new_n_n829_ = new_n_n350_ & new_n_n432_ & new_n_n82_;
  assign new_na8_ = new_n_n408_ & new_no0_ & new_n_n91_;
  assign new_nd8_ = new_n_n408_ & new_no0_ & new_n_n94_;
  assign new_nk8_ = new_n_n820_ | new_n_n821_;
  assign new_n_n814_ = new_no0_ & new_n_n112_ & new_n_n147_;
  assign new_n_n807_ = new_n_n194_ & new_n_n119_ & new_n_n145_;
  assign new_n_n774_ = new_n_n157_ & new_nz3_;
  assign new_nn9_ = new_n_n411_ | new_n_n170_ | new_n_n767_;
  assign new_ny15_ = new_nq0_ | new_n_n411_ | new_n_n199_;
  assign new_ny17_ = new_n_n732_ | new_n_n742_ | new_n_n697_;
  assign new_n_n728_ = new_nm0_ & new_no0_ & new_n_n408_;
  assign new_n_n652_ = new_n_n281_ & new_n_n283_ & new_n_n282_;
  assign new_n_n648_ = new_nl0_ & new_n_n431_;
  assign new_na24_ = new_n_n639_ | new_n_n640_;
  assign new_n_n633_ = new_n_n365_ & new_nu2_ & new_n_n306_;
  assign new_n_n613_ = new_n_n302_ & new_na17_ & new_n_n303_;
  assign new_nn25_ = new_nj6_ & new_ni6_ & new_nh6_;
  assign new_n_n592_ = new_nl1_ & new_nk1_;
  assign new_nj26_ = new_nq0_ | new_n_n422_;
  assign new_na27_ = new_n_n439_ | new_n_n320_ | new_nj25_;
  assign new_n_n586_ = new_n_n327_ & new_n_n396_;
  assign new_np28_ = new_n_n579_ | new_n_n333_;
  assign new_n_n566_ = new_nn0_ & new_n_n408_ & new_n_n341_;
  assign new_n_n563_ = new_n_n346_ & new_n_n441_ & new_n_n348_;
  assign new_nq29_ = new_nx3_ | new_na17_ | new_n_n351_;
  assign new_nv29_ = new_n_n365_ | new_n_n437_ | new_n_n458_;
  assign new_nb31_ = new_n_n404_ & new_nl25_ & new_n_n368_;
  assign new_nl31_ = new_n_n439_ | new_nf4_ | new_n_n461_;
  assign new_n_n540_ = new_n_n431_ & new_nl0_ & new_nm0_;
  assign new_ni32_ = new_n_n537_ | new_n_n386_;
  assign new_n_n532_ = new_n_n392_ & new_n_n391_ & new_n_n390_;
  assign new_nt32_ = new_nj6_ & new_nt0_ & new_n_n401_;
  assign new_nd33_ = new_n_n449_ | new_n_n409_ | new_n_n523_;
  assign new_n_n505_ = new_n_n425_ & new_nl0_;
  assign new_n_n498_ = new_n_n431_ & new_n_n430_ & new_n_n422_;
  assign new_n_n491_ = new_nk0_ & new_nl0_ & new_n_n426_;
  assign new_ne34_ = new_n_n439_ & new_nk1_ & new_n_n432_;
  assign new_nh34_ = new_n_n484_ | new_n_n485_;
  assign new_nr34_ = new_nj1_ & new_nl4_;
  assign new_n_n478_ = new_nj6_ & new_na1_ & new_nl6_;
  assign new_ne35_ = new_n_n445_ | new_nh4_;
  assign new_n_n453_ = ~new_nl35_;
  assign new_n_n444_ = ~new_na1_;
  assign new_n_n435_ = ~new_nf1_;
  assign new_n_n424_ = ~new_nh3_;
  assign new_n_n421_ = ~new_ne3_;
  assign new_n_n410_ = ~new_nx0_;
  assign new_n_n400_ = ~new_nu0_;
  assign new_n_n389_ = ~new_no32_;
  assign new_n_n360_ = ~new_nd30_;
  assign new_n_n349_ = ~new_nq29_;
  assign new_n_n338_ = ~new_no25_;
  assign new_n_n327_ = ~new_ns28_;
  assign new_n_n324_ = ~new_nu3_;
  assign new_n_n313_ = ~new_nk25_;
  assign new_n_n302_ = ~new_ny2_;
  assign new_n_n291_ = ~new_nd24_;
  assign new_n_n275_ = ~new_na23_;
  assign new_n_n261_ = ~new_ns21_;
  assign new_n_n250_ = ~new_na21_;
  assign new_n_n239_ = ~new_nc2_;
  assign new_n_n228_ = ~new_nx18_;
  assign new_n_n214_ = ~new_no17_;
  assign new_n_n203_ = ~new_nm16_;
  assign new_n_n192_ = ~new_ne33_;
  assign new_n_n176_ = ~new_nn31_;
  assign new_n_n165_ = ~new_nl30_;
  assign new_n_n162_ = ~new_nm30_;
  assign new_n_n151_ = ~new_nl28_;
  assign new_n_n140_ = ~new_nw27_;
  assign new_n_n129_ = ~new_ng27_;
  assign new_n_n104_ = ~new_nd25_;
  assign new_n_n93_ = ~new_ny23_;
  assign new_n_n1_ = ~new_ni33_;
  assign new_n_n1104_ = new_n_n0_ & new_n_n428_;
  assign new_n_n1064_ = new_nn1_ & new_n_n356_;
  assign new_n_n1043_ = new_n_n30_ & new_n_n32_ & new_n_n29_;
  assign new_n_n1036_ = new_n_n35_ & new_n_n34_;
  assign new_n_n1025_ = new_n_n37_ & new_n_n83_ & new_n_n38_;
  assign new_n_n1017_ = new_na17_ & new_n_n83_ & new_n_n40_;
  assign new_n_n990_ = new_na17_ & new_n_n83_ & new_n_n46_;
  assign new_n_n982_ = new_n_n350_ & new_n_n432_ & new_n_n48_;
  assign new_n_n970_ = new_n_n350_ & new_n_n83_ & new_n_n50_;
  assign new_n_n962_ = new_n_n51_ & new_n_n83_ & new_n_n52_;
  assign new_n_n958_ = new_n_n350_ & new_nv1_ & new_n_n54_;
  assign new_n_n950_ = new_n_n55_ & new_nw1_ & new_n_n56_;
  assign new_n_n938_ = new_n_n57_ & new_n_n432_ & new_n_n58_;
  assign new_n_n930_ = new_na17_ & new_n_n432_ & new_n_n60_;
  assign new_n_n907_ = new_n_n350_ & new_n_n83_ & new_n_n64_;
  assign new_n_n903_ = new_na17_ & new_n_n432_ & new_n_n66_;
  assign new_n_n895_ = new_n_n350_ & new_nc2_ & new_n_n68_;
  assign new_n_n883_ = new_n_n350_ & new_n_n432_ & new_n_n70_;
  assign new_n_n875_ = new_n_n71_ & new_n_n432_ & new_n_n72_;
  assign new_no7_ = new_n_n869_ | new_n_n867_ | new_n_n866_ | new_n_n868_ | new_n_n870_ | new_n_n865_ | new_n_n864_ | new_n_n863_ | new_n_n862_;
  assign new_n_n851_ = new_n_n77_ & new_nh2_ & new_n_n78_;
  assign new_n_n843_ = new_na17_ & new_ni2_ & new_n_n80_;
  assign new_n_n828_ = new_na17_ & new_n_n83_ & new_n_n82_;
  assign new_nz7_ = new_n_n408_ & new_no0_ & new_n_n90_;
  assign new_ne8_ = new_n_n408_ & new_no0_ & new_n_n95_;
  assign new_n_n822_ = new_no0_ & new_n_n104_ & new_n_n147_;
  assign new_no8_ = new_n_n812_ | new_n_n813_;
  assign new_nr8_ = new_n_n806_ | new_n_n807_;
  assign new_nj9_ = new_n_n408_ & new_no0_ & new_n_n158_;
  assign new_n_n768_ = new_n_n432_ & new_no0_ & new_n_n169_;
  assign new_nk15_ = new_n_n378_ | new_ne1_ | new_nd1_;
  assign new_n_n732_ = new_ne0_ & new_no0_ & new_n_n408_;
  assign new_ni18_ = new_n_n728_ | new_n_n742_ | new_n_n697_;
  assign new_n_n651_ = new_n_n387_ & new_n_n283_ & new_n_n282_;
  assign new_nu23_ = new_n_n378_ | new_n_n648_ | new_n_n647_;
  assign new_n_n640_ = new_nj_ & new_n_n305_ & new_n_n353_;
  assign new_n_n634_ = new_nk_ & new_n_n305_ & new_n_n353_;
  assign new_nz24_ = new_n_n608_ | new_nw16_;
  assign new_no25_ = new_nk6_ & new_nl6_;
  assign new_n_n593_ = new_nl1_ & new_nj1_;
  assign new_nl26_ = new_n_n439_ | new_n_n424_ | new_nj25_;
  assign new_ny26_ = new_nq0_ | new_n_n427_;
  assign new_nk28_ = new_nq0_ | new_n_n328_;
  assign new_n_n580_ = new_nk6_ & new_nl25_ & new_n_n332_;
  assign new_nf29_ = new_n_n342_ & new_nl4_;
  assign new_nn29_ = new_n_n562_ | new_n_n560_ | new_n_n559_ | new_n_n561_ | new_n_n563_ | new_n_n558_ | new_n_n557_ | new_n_n556_ | new_n_n555_;
  assign new_nr29_ = new_n_n553_ | new_n_n551_ | new_n_n550_ | new_n_n552_ | new_n_n554_;
  assign new_nu29_ = new_na17_ | new_nx3_;
  assign new_nc31_ = new_n_n408_ & new_no4_ & new_n_n369_;
  assign new_nk31_ = new_nj25_ | new_nd4_;
  assign new_nc32_ = new_n_n439_ | new_ng4_ | new_n_n460_;
  assign new_n_n537_ = new_nn1_ & new_ni4_;
  assign new_n_n533_ = new_n_n389_ & new_n_n391_ & new_n_n390_;
  assign new_nu32_ = new_nn4_ & new_nk4_ & new_n_n402_;
  assign new_nc33_ = new_na17_ | new_nq0_ | new_n_n411_;
  assign new_nr33_ = new_n_n504_ | new_n_n503_ | new_n_n502_;
  assign new_n_n499_ = new_nk0_ & new_nl0_ & new_n_n422_;
  assign new_n_n490_ = new_n_n431_ & new_n_n430_ & new_n_n426_;
  assign new_nd34_ = new_n_n439_ & new_nj1_ & new_n_n432_;
  assign new_n_n485_ = new_ni4_ & new_n_n435_;
  assign new_nq34_ = new_ni1_ & new_nl4_;
  assign new_n_n477_ = new_nz0_ & new_nk6_ & new_nl6_;
  assign new_n_n470_ = new_n_n452_ & new_nl1_;
  assign new_n_n452_ = ~new_nb1_;
  assign new_n_n445_ = ~new_nf35_;
  assign new_n_n434_ = ~new_nc4_;
  assign new_n_n425_ = ~new_ni3_;
  assign new_n_n420_ = ~new_nq3_;
  assign new_n_n411_ = ~new_no0_;
  assign new_n_n399_ = ~new_ns32_;
  assign new_n_n390_ = ~new_nr32_;
  assign new_n_n359_ = ~new_ne30_;
  assign new_n_n350_ = ~new_ns16_;
  assign new_n_n337_ = ~new_nv28_;
  assign new_n_n328_ = ~new_nw3_;
  assign new_n_n323_ = ~new_np3_;
  assign new_n_n314_ = ~new_nr35_;
  assign new_n_n301_ = ~new_np23_;
  assign new_n_n292_ = ~new_nv2_;
  assign new_n_n265_ = ~new_nh22_;
  assign new_n_n260_ = ~new_nr21_;
  assign new_n_n251_ = ~new_ni2_;
  assign new_n_n238_ = ~new_nw19_;
  assign new_n_n229_ = ~new_nx1_;
  assign new_n_n224_ = ~new_nn18_;
  assign new_n_n202_ = ~new_nh16_;
  assign new_n_n193_ = ~new_nd33_;
  assign new_n_n175_ = ~new_no31_;
  assign new_n_n166_ = ~new_nk30_;
  assign new_n_n161_ = ~new_na30_;
  assign new_n_n152_ = ~new_nk28_;
  assign new_n_n139_ = ~new_nv27_;
  assign new_n_n130_ = ~new_nh27_;
  assign new_n_n103_ = ~new_nb25_;
  assign new_n_n94_ = ~new_nc24_;
  assign new_n_n2_ = ~new_nh33_;
  assign new_n_n1096_ = new_n_n6_ & new_n_n428_;
  assign new_n_n1087_ = new_nk0_ & new_nl0_ & new_n_n12_;
  assign new_np6_ = new_n_n206_ & new_n_n408_ & new_no0_;
  assign new_nt6_ = new_n_n1041_ | new_n_n1039_ | new_n_n1038_ | new_n_n1037_ | new_n_n1040_ | new_n_n1042_;
  assign new_n_n1034_ = new_n_n36_ & new_nm1_;
  assign new_n_n1028_ = new_n_n37_ & new_n_n432_ & new_n_n38_;
  assign new_n_n1018_ = new_n_n350_ & new_n_n432_ & new_n_n40_;
  assign new_n_n989_ = new_n_n45_ & new_n_n83_ & new_n_n46_;
  assign new_n_n979_ = new_n_n350_ & new_n_n83_ & new_n_n48_;
  assign new_n_n973_ = new_n_n350_ & new_n_n432_ & new_n_n50_;
  assign new_n_n963_ = new_na17_ & new_n_n83_ & new_n_n52_;
  assign new_n_n957_ = new_na17_ & new_n_n432_ & new_n_n54_;
  assign new_n_n947_ = new_n_n55_ & new_n_n432_ & new_n_n56_;
  assign new_n_n941_ = new_n_n57_ & new_nx1_ & new_n_n58_;
  assign new_n_n931_ = new_n_n350_ & new_ny1_ & new_n_n60_;
  assign new_n_n918_ = new_na17_ & new_n_n83_ & new_n_n62_;
  assign new_n_n908_ = new_n_n63_ & new_n_n83_ & new_n_n64_;
  assign new_n_n902_ = new_n_n65_ & new_n_n432_ & new_n_n66_;
  assign new_n_n892_ = new_n_n350_ & new_n_n432_ & new_n_n68_;
  assign new_n_n886_ = new_n_n350_ & new_nd2_ & new_n_n70_;
  assign new_n_n876_ = new_na17_ & new_n_n432_ & new_n_n72_;
  assign new_n_n870_ = new_na17_ & new_nf2_ & new_n_n74_;
  assign new_n_n860_ = new_n_n75_ & new_ng2_ & new_n_n76_;
  assign new_nr7_ = new_n_n842_ | new_n_n840_ | new_n_n839_ | new_n_n841_ | new_n_n843_ | new_n_n838_ | new_n_n837_ | new_n_n836_ | new_n_n835_;
  assign new_n_n831_ = new_na17_ & new_n_n432_ & new_n_n82_;
  assign new_ny7_ = new_n_n408_ & new_no0_ & new_n_n89_;
  assign new_nf8_ = new_n_n408_ & new_no0_ & new_n_n96_;
  assign new_n_n820_ = new_no0_ & new_n_n106_ & new_n_n147_;
  assign new_nn8_ = new_n_n814_ | new_n_n815_;
  assign new_n_n808_ = new_no0_ & new_n_n118_ & new_n_n147_;
  assign new_n_n775_ = new_n_n155_ & new_ny3_;
  assign new_n_n769_ = new_no0_ & new_n_n168_ & new_n_n167_;
  assign new_nt9_ = new_n_n434_ & new_n_n433_ & new_n_n190_;
  assign new_no23_ = new_nt2_ & new_nl4_;
  assign new_nw23_ = new_n_n645_ | new_n_n646_;
  assign new_n_n641_ = new_n_n387_ & new_n_n288_ & new_n_n287_;
  assign new_ne24_ = new_n_n633_ | new_n_n634_;
  assign new_n_n605_ = new_nh6_ & new_ni6_ & new_n_n311_;
  assign new_np25_ = new_nj6_ & new_ni6_ & new_n_n401_;
  assign new_nw25_ = new_n_n439_ | new_n_n415_ | new_nj25_;
  assign new_ng26_ = new_nq0_ | new_n_n421_;
  assign new_nx26_ = new_n_n439_ | new_n_n429_ | new_nj25_;
  assign new_n_n575_ = new_n_n400_ & new_nj1_ & new_n_n336_;
  assign new_n_n568_ = new_nl4_ & new_nx3_ & new_n_n387_;
  assign new_ng29_ = new_ny3_ | new_nx3_ | new_na17_;
  assign new_n_n561_ = new_n_n350_ & new_n_n441_ & new_n_n348_;
  assign new_no29_ = new_ny3_ & new_n_n440_ & new_n_n387_;
  assign new_n_n548_ = new_n_n378_ & new_n_n355_ & new_n_n354_;
  assign new_nd31_ = new_n_n543_ | new_nz29_;
  assign new_ns31_ = new_n_n380_ & new_no0_;
  assign new_nb32_ = new_n_n461_ | new_nd4_ | new_nj25_;
  assign new_nj32_ = new_n_n387_ & new_n_n408_ & new_no0_;
  assign new_np32_ = new_n_n531_ | new_n_n530_ | new_n_n529_;
  assign new_n_n527_ = new_nh6_ & new_n_n400_ & new_n_n399_;
  assign new_nb33_ = new_n_n408_ & new_nm1_;
  assign new_n_n504_ = new_n_n419_ & new_nl0_;
  assign new_n_n497_ = new_nk0_ & new_nl0_ & new_n_n423_;
  assign new_n_n492_ = new_n_n431_ & new_n_n430_ & new_n_n425_;
  assign new_nc34_ = new_n_n439_ & new_ni1_ & new_n_n432_;
  assign new_n_n484_ = new_n_n436_ & new_nf1_;
  assign new_nt34_ = new_nl1_ & new_nl4_;
  assign new_n_n480_ = new_nj6_ & new_nk6_ & new_nb1_;
  assign new_n_n471_ = new_n_n444_ & new_nk1_;
  assign new_nk35_ = new_n_n457_ & new_n_n456_ & new_n_n453_;
  assign new_n_n451_ = ~new_nk35_;
  assign new_n_n442_ = ~new_nd35_;
  assign new_n_n437_ = ~new_nz3_;
  assign new_n_n426_ = ~new_nj3_;
  assign new_n_n419_ = ~new_na3_;
  assign new_n_n408_ = ~new_nq0_;
  assign new_n_n401_ = ~new_nt25_;
  assign new_n_n391_ = ~new_nq32_;
  assign new_n_n376_ = ~new_nu31_;
  assign new_n_n365_ = ~new_nl4_;
  assign new_n_n358_ = ~new_nf30_;
  assign new_n_n347_ = ~new_np29_;
  assign new_n_n340_ = ~new_nb29_;
  assign new_n_n329_ = ~new_nm28_;
  assign new_n_n322_ = ~new_no3_;
  assign new_n_n311_ = ~new_nh25_;
  assign new_n_n304_ = ~new_nt24_;
  assign new_n_n293_ = ~new_ni24_;
  assign new_n_n277_ = ~new_nj23_;
  assign new_n_n266_ = ~new_nf22_;
  assign new_n_n259_ = ~new_nt21_;
  assign new_n_n248_ = ~new_nv20_;
  assign new_n_n241_ = ~new_nd2_;
  assign new_n_n230_ = ~new_nc19_;
  assign new_n_n223_ = ~new_nu1_;
  assign new_n_n212_ = ~new_nj17_;
  assign new_n_n194_ = ~new_na25_;
  assign new_n_n178_ = ~new_np31_;
  assign new_n_n167_ = ~new_nu30_;
  assign new_n_n160_ = ~new_nb30_;
  assign new_n_n149_ = ~new_ni28_;
  assign new_n_n142_ = ~new_nz27_;
  assign new_n_n131_ = ~new_nj27_;
  assign new_n_n124_ = ~new_ny26_;
  assign new_n_n113_ = ~new_ni26_;
  assign new_n_n3_ = ~new_nm33_;
  assign new_n_n1095_ = new_n_n431_ & new_n_n8_ & new_n_n6_;
  assign new_n_n1088_ = new_n_n12_ & new_nm3_;
  assign new_n_n1049_ = new_n_n28_ & new_n_n32_ & new_n_n27_;
  assign new_n_n1042_ = new_n_n378_ & new_no4_ & new_n_n31_;
  assign new_nv6_ = new_n_n1033_ | new_n_n1034_;
  assign new_n_n1027_ = new_n_n350_ & new_n_n432_ & new_n_n38_;
  assign new_n_n1019_ = new_n_n39_ & new_n_n432_ & new_n_n40_;
  assign new_n_n988_ = new_n_n350_ & new_n_n83_ & new_n_n46_;
  assign new_n_n980_ = new_n_n47_ & new_n_n83_ & new_n_n48_;
  assign new_n_n972_ = new_na17_ & new_n_n83_ & new_n_n50_;
  assign new_n_n964_ = new_n_n350_ & new_n_n432_ & new_n_n52_;
  assign new_n_n956_ = new_n_n53_ & new_n_n432_ & new_n_n54_;
  assign new_n_n948_ = new_na17_ & new_n_n432_ & new_n_n56_;
  assign new_n_n940_ = new_n_n350_ & new_nx1_ & new_n_n58_;
  assign new_n_n932_ = new_n_n59_ & new_ny1_ & new_n_n60_;
  assign new_n_n917_ = new_n_n61_ & new_n_n83_ & new_n_n62_;
  assign new_n_n909_ = new_na17_ & new_n_n83_ & new_n_n64_;
  assign new_n_n901_ = new_n_n350_ & new_n_n432_ & new_n_n66_;
  assign new_n_n893_ = new_n_n67_ & new_n_n432_ & new_n_n68_;
  assign new_n_n885_ = new_na17_ & new_n_n432_ & new_n_n70_;
  assign new_n_n877_ = new_n_n350_ & new_ne2_ & new_n_n72_;
  assign new_n_n869_ = new_n_n73_ & new_nf2_ & new_n_n74_;
  assign new_n_n861_ = new_na17_ & new_ng2_ & new_n_n76_;
  assign new_nq7_ = new_n_n851_ | new_n_n849_ | new_n_n848_ | new_n_n850_ | new_n_n852_ | new_n_n847_ | new_n_n846_ | new_n_n845_ | new_n_n844_;
  assign new_n_n830_ = new_n_n81_ & new_n_n432_ & new_n_n82_;
  assign new_nx7_ = new_n_n408_ & new_no0_ & new_n_n88_;
  assign new_ng8_ = new_n_n408_ & new_no0_ & new_n_n97_;
  assign new_n_n821_ = new_n_n194_ & new_n_n105_ & new_n_n145_;
  assign new_n_n815_ = new_n_n194_ & new_n_n111_ & new_n_n145_;
  assign new_n_n809_ = new_n_n194_ & new_n_n117_ & new_n_n145_;
  assign new_ni9_ = new_n_n411_ | new_n_n156_ | new_n_n774_;
  assign new_nm9_ = new_n_n768_ | new_n_n769_;
  assign new_n_n764_ = new_no0_ & new_n_n178_ & new_n_n177_;
  assign new_np23_ = new_nn0_ | new_nm0_ | new_n_n284_;
  assign new_n_n647_ = new_n_n430_ & new_nk0_;
  assign new_nz23_ = new_nu2_ & new_nl4_;
  assign new_nd24_ = new_nv2_ & new_nl4_;
  assign new_nj25_ = new_n_n314_ & new_n_n457_;
  assign new_nq25_ = new_nl6_ & new_nk6_ & new_nj6_;
  assign new_nt25_ = new_nk1_ | new_nl1_;
  assign new_ni26_ = new_n_n439_ | new_n_n423_ | new_nj25_;
  assign new_nv26_ = new_nq0_ | new_n_n426_;
  assign new_n_n574_ = new_n_n393_ & new_nj6_ & new_n_n336_;
  assign new_na29_ = new_n_n568_ | new_n_n340_;
  assign new_ni29_ = new_n_n440_ & new_n_n387_ & new_n_n343_;
  assign new_n_n562_ = new_n_n347_ & new_n_n441_ & new_n_n348_;
  assign new_np29_ = new_nl4_ & new_n_n441_ & new_nz3_;
  assign new_n_n549_ = new_nn0_ & new_nt15_;
  assign new_nm31_ = new_n_n439_ | new_n_n461_ | new_nd4_;
  assign new_nt31_ = new_nn0_ | new_n_n540_ | new_n_n539_;
  assign new_n_n538_ = new_nl25_ & new_n_n385_ & new_n_n384_;
  assign new_nk32_ = new_nq0_ | new_n_n411_ | new_n_n388_;
  assign new_no32_ = new_ni6_ & new_nj6_;
  assign new_ns32_ = new_nl1_ | new_nk1_ | new_ni1_;
  assign new_na33_ = new_n_n411_ | new_n_n406_ | new_n_n407_;
  assign new_n_n503_ = new_n_n425_ & new_n_n430_;
  assign new_nv33_ = new_n_n428_ | new_n_n497_ | new_n_n496_;
  assign new_ny33_ = new_n_n428_ | new_n_n491_ | new_n_n490_;
  assign new_nb34_ = new_n_n439_ & new_nh1_ & new_n_n432_;
  assign new_ni34_ = new_n_n437_ | new_n_n458_ | new_n_n438_;
  assign new_ns34_ = new_nk1_ & new_nl4_;
  assign new_n_n479_ = new_nz0_ & new_na1_ & new_nl6_;
  assign new_nd35_ = new_n_n443_ | new_n_n471_ | new_n_n470_;
  assign new_n_n459_ = ~new_nw34_;
  assign new_n_n450_ = ~new_ni35_;
  assign new_n_n443_ = ~new_ne35_;
  assign new_n_n436_ = ~new_ni4_;
  assign new_n_n427_ = ~new_nk3_;
  assign new_n_n418_ = ~new_nr3_;
  assign new_n_n409_ = ~new_nb35_;
  assign new_nh6_ = ~new_nh1_;
  assign new_n_n392_ = ~new_np32_;
  assign new_n_n375_ = ~new_nw31_;
  assign new_n_n366_ = ~new_nx30_;
  assign new_n_n357_ = ~new_nh30_;
  assign new_n_n348_ = ~new_nr29_;
  assign new_n_n339_ = ~new_nx28_;
  assign new_n_n330_ = ~new_nf25_;
  assign new_n_n321_ = ~new_nn3_;
  assign new_n_n312_ = ~new_ni25_;
  assign new_n_n303_ = ~new_nu24_;
  assign new_n_n294_ = ~new_nh24_;
  assign new_n_n276_ = ~new_nb23_;
  assign new_n_n267_ = ~new_ng22_;
  assign new_n_n258_ = ~new_nj21_;
  assign new_n_n249_ = ~new_nh2_;
  assign new_n_n240_ = ~new_nb20_;
  assign new_n_n231_ = ~new_ny1_;
  assign new_n_n222_ = ~new_ni18_;
  assign new_n_n213_ = ~new_np1_;
  assign new_n_n204_ = ~new_ne1_;
  assign new_n_n177_ = ~new_nq31_;
  assign new_n_n168_ = ~new_nt30_;
  assign new_n_n159_ = ~new_nx29_;
  assign new_n_n150_ = ~new_nh28_;
  assign new_n_n141_ = ~new_ny27_;
  assign new_n_n132_ = ~new_nk27_;
  assign new_n_n123_ = ~new_nx26_;
  assign new_n_n114_ = ~new_nj26_;
  assign new_n_n4_ = ~new_nl33_;
  assign new_n_n1097_ = new_n_n5_ & new_n_n4_ & new_n_n3_;
  assign new_nv4_ = new_n_n1088_ | new_n_n1087_ | new_n_n1086_;
  assign new_nq6_ = new_n_n1055_ | new_n_n1056_;
  assign new_n_n1048_ = new_n_n378_ & new_no4_ & new_n_n29_;
  assign new_n_n1038_ = new_nn0_ & new_n_n32_ & new_n_n31_;
  assign new_n_n1030_ = new_n_n350_ & new_nn1_ & new_n_n38_;
  assign new_n_n1020_ = new_na17_ & new_n_n432_ & new_n_n40_;
  assign new_ng7_ = new_n_n941_ | new_n_n939_ | new_n_n938_ | new_n_n940_ | new_n_n942_ | new_n_n937_ | new_n_n936_ | new_n_n935_ | new_n_n934_;
  assign new_n_n933_ = new_na17_ & new_ny1_ & new_n_n60_;
  assign new_n_n79_ = ~new_nx20_;
  assign new_n_n68_ = ~new_nv19_;
  assign new_n_n57_ = ~new_nu18_;
  assign new_n_n46_ = ~new_ns17_;
  assign new_n_n35_ = ~new_nl16_;
  assign new_nr4_ = new_n_n1093_ | new_n_n1095_ | new_n_n1094_ | new_n_n1096_;
  assign new_n_n1089_ = new_n_n11_ & new_n_n10_ & new_n_n9_;
  assign new_n_n1063_ = new_nn1_ & new_n_n438_;
  assign new_n_n1047_ = new_nn0_ & new_no4_ & new_n_n29_;
  assign new_n_n1039_ = new_n_n378_ & new_n_n32_ & new_n_n31_;
  assign new_n_n1029_ = new_na17_ & new_n_n432_ & new_n_n38_;
  assign new_n_n1021_ = new_n_n350_ & new_no1_ & new_n_n40_;
  assign new_n_n942_ = new_na17_ & new_nx1_ & new_n_n58_;
  assign new_nh7_ = new_n_n932_ | new_n_n930_ | new_n_n929_ | new_n_n931_ | new_n_n933_ | new_n_n928_ | new_n_n927_ | new_n_n926_ | new_n_n925_;
  assign new_n_n80_ = ~new_nz20_;
  assign new_n_n67_ = ~new_nt19_;
  assign new_n_n58_ = ~new_nw18_;
  assign new_n_n45_ = ~new_nq17_;
  assign new_n_n36_ = ~new_np16_;
  assign new_np4_ = new_n_n1101_ | new_n_n1103_ | new_n_n1102_ | new_n_n1104_;
  assign new_n_n1099_ = new_n_n431_ & new_n_n5_ & new_n_n3_;
  assign new_n_n1090_ = new_nk0_ & new_n_n10_ & new_n_n9_;
  assign new_ne5_ = new_nm0_ & new_nn3_;
  assign new_n_n1046_ = new_n_n30_ & new_no4_ & new_n_n29_;
  assign new_nu6_ = new_n_n1035_ | new_n_n1036_;
  assign new_n_n1032_ = new_na17_ & new_nn1_ & new_n_n38_;
  assign new_n_n1022_ = new_n_n39_ & new_no1_ & new_n_n40_;
  assign new_ne7_ = new_n_n959_ | new_n_n957_ | new_n_n956_ | new_n_n958_ | new_n_n960_ | new_n_n955_ | new_n_n954_ | new_n_n953_ | new_n_n952_;
  assign new_n_n951_ = new_na17_ & new_nw1_ & new_n_n56_;
  assign new_n_n81_ = ~new_nc21_;
  assign new_n_n66_ = ~new_nq19_;
  assign new_n_n55_ = ~new_np18_;
  assign new_n_n48_ = ~new_nx17_;
  assign new_n_n37_ = ~new_nr16_;
  assign new_n_n1098_ = new_nk0_ & new_n_n4_ & new_n_n3_;
  assign new_n_n1091_ = new_n_n431_ & new_n_n11_ & new_n_n9_;
  assign new_n_n1071_ = new_n_n431_ & new_n_n430_ & new_n_n17_;
  assign new_n_n1045_ = new_n_n378_ & new_n_n32_ & new_n_n29_;
  assign new_n_n1037_ = new_n_n33_ & new_n_n32_ & new_n_n31_;
  assign new_n_n1031_ = new_n_n37_ & new_nn1_ & new_n_n38_;
  assign new_n_n1023_ = new_na17_ & new_no1_ & new_n_n40_;
  assign new_n_n960_ = new_na17_ & new_nv1_ & new_n_n54_;
  assign new_nf7_ = new_n_n950_ | new_n_n948_ | new_n_n947_ | new_n_n949_ | new_n_n951_ | new_n_n946_ | new_n_n945_ | new_n_n944_ | new_n_n943_;
  assign new_n_n82_ = ~new_ne21_;
  assign new_n_n65_ = ~new_no19_;
  assign new_n_n56_ = ~new_nr18_;
  assign new_n_n47_ = ~new_nv17_;
  assign new_n_n38_ = ~new_nv16_;
  assign new_n_n0_ = ~new_nj33_;
  assign new_nq4_ = new_n_n1097_ | new_n_n1099_ | new_n_n1098_ | new_n_n1100_;
  assign new_n_n1092_ = new_n_n9_ & new_n_n428_;
  assign new_nb5_ = new_n_n1070_ | new_n_n1069_ | new_n_n1068_;
  assign new_ng5_ = new_nm0_ & new_np3_;
  assign new_n_n1060_ = new_n_n20_ & new_n_n438_;
  assign new_n_n1054_ = new_n_n378_ & new_no4_ & new_n_n27_;
  assign new_nx6_ = new_n_n1022_ | new_n_n1020_ | new_n_n1019_ | new_n_n1021_ | new_n_n1023_ | new_n_n1018_ | new_n_n1017_ | new_n_n1016_ | new_n_n1015_;
  assign new_nc7_ = new_n_n977_ | new_n_n975_ | new_n_n974_ | new_n_n976_ | new_n_n978_ | new_n_n973_ | new_n_n972_ | new_n_n971_ | new_n_n970_;
  assign new_n_n969_ = new_na17_ & new_nu1_ & new_n_n52_;
  assign new_nh18_ = new_n_n729_ | new_n_n222_;
  assign new_n_n725_ = new_n_n227_ & new_n_n378_ & new_n_n254_;
  assign new_n_n646_ = new_nk0_ & new_nl0_ & new_nt15_;
  assign new_nc24_ = new_n_n635_ | new_n_n637_ | new_n_n636_ | new_n_n638_;
  assign new_no26_ = new_n_n439_ | new_n_n425_ | new_nj25_;
  assign new_n_n83_ = ~new_nu16_;
  assign new_n_n28_ = ~new_nw15_;
  assign new_nc6_ = ~new_np34_;
  assign new_no5_ = ~new_nc34_;
  assign new_n_n10_ = ~new_nr33_;
  assign new_n_n1100_ = new_n_n3_ & new_n_n428_;
  assign new_ns4_ = new_n_n1089_ | new_n_n1091_ | new_n_n1090_ | new_n_n1092_;
  assign new_n_n1070_ = new_n_n18_ & new_ns3_;
  assign new_nf5_ = new_nm0_ & new_no3_;
  assign new_n_n1059_ = new_n_n20_ & new_n_n21_;
  assign new_nr6_ = new_n_n1053_ | new_n_n1051_ | new_n_n1050_ | new_n_n1049_ | new_n_n1052_ | new_n_n1054_;
  assign new_nw6_ = new_n_n1031_ | new_n_n1029_ | new_n_n1028_ | new_n_n1030_ | new_n_n1032_ | new_n_n1027_ | new_n_n1026_ | new_n_n1025_ | new_n_n1024_;
  assign new_n_n978_ = new_na17_ & new_nt1_ & new_n_n50_;
  assign new_nd7_ = new_n_n968_ | new_n_n966_ | new_n_n965_ | new_n_n967_ | new_n_n969_ | new_n_n964_ | new_n_n963_ | new_n_n962_ | new_n_n961_;
  assign new_n_n729_ = new_n_n223_ & new_n_n378_ & new_n_n254_;
  assign new_nr18_ = new_n_n725_ | new_n_n226_;
  assign new_n_n645_ = new_n_n431_ & new_n_n430_ & new_nt15_;
  assign new_n_n639_ = new_n_n365_ & new_nt2_ & new_n_n306_;
  assign new_nz25_ = new_n_n439_ | new_n_n413_ | new_nj25_;
  assign new_n_n84_ = ~new_nh21_;
  assign new_n_n27_ = ~new_ny15_;
  assign new_nd6_ = ~new_nq34_;
  assign new_nn5_ = ~new_nb34_;
  assign new_n_n11_ = ~new_nq33_;
  assign new_n_n1102_ = new_nk0_ & new_n_n1_ & new_n_n0_;
  assign new_n_n1093_ = new_n_n8_ & new_n_n7_ & new_n_n6_;
  assign new_n_n1069_ = new_nk0_ & new_nl0_ & new_n_n18_;
  assign new_ni5_ = new_nm0_ & new_nr3_;
  assign new_n_n1062_ = new_nn1_ & new_n_n21_;
  assign new_n_n1055_ = new_no0_ & new_n_n26_ & new_n_n25_;
  assign new_n_n1040_ = new_n_n33_ & new_no4_ & new_n_n31_;
  assign new_na7_ = new_n_n995_ | new_n_n993_ | new_n_n992_ | new_n_n994_ | new_n_n996_ | new_n_n991_ | new_n_n990_ | new_n_n989_ | new_n_n988_;
  assign new_n_n987_ = new_na17_ & new_ns1_ & new_n_n48_;
  assign new_n_n771_ = new_n_n164_ & new_n_n163_ & new_n_n180_;
  assign new_n_n730_ = new_nd0_ & new_no0_ & new_n_n408_;
  assign new_np18_ = new_n_n229_ & new_nl4_;
  assign new_nj23_ = new_nr2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n650_ = new_ni_ & new_n_n305_ & new_n_n353_;
  assign new_n_n597_ = new_n_n319_ & new_ni1_;
  assign new_n_n26_ = ~new_nl15_;
  assign new_na6_ = ~new_nn34_;
  assign new_nq5_ = ~new_ne34_;
  assign new_n_n12_ = ~new_nt33_;
  assign new_n_n1101_ = new_n_n2_ & new_n_n1_ & new_n_n0_;
  assign new_n_n1094_ = new_nk0_ & new_n_n7_ & new_n_n6_;
  assign new_n_n1068_ = new_n_n431_ & new_n_n430_ & new_n_n18_;
  assign new_nh5_ = new_nm0_ & new_nq3_;
  assign new_n_n1061_ = new_n_n20_ & new_n_n356_;
  assign new_n_n1056_ = new_n_n432_ & new_n_n24_ & new_n_n23_;
  assign new_ns6_ = new_n_n1047_ | new_n_n1045_ | new_n_n1044_ | new_n_n1043_ | new_n_n1046_ | new_n_n1048_;
  assign new_n_n996_ = new_na17_ & new_nr1_ & new_n_n46_;
  assign new_nb7_ = new_n_n986_ | new_n_n984_ | new_n_n983_ | new_n_n985_ | new_n_n987_ | new_n_n982_ | new_n_n981_ | new_n_n980_ | new_n_n979_;
  assign new_n_n765_ = new_n_n176_ & new_n_n175_ & new_n_n180_;
  assign new_nf18_ = new_n_n225_ & new_nl4_;
  assign new_n_n726_ = new_nk0_ & new_no0_ & new_n_n408_;
  assign new_n_n656_ = new_nl4_ & new_n_n387_;
  assign new_nq23_ = new_n_n649_ | new_n_n650_;
  assign new_nk25_ = new_n_n412_ | new_n_n315_ | new_n_n599_;
  assign new_n_n25_ = ~new_nm15_;
  assign new_nb6_ = ~new_no34_;
  assign new_np5_ = ~new_nd34_;
  assign new_n_n13_ = ~new_nu33_;
  assign new_n_n1084_ = new_nk0_ & new_nl0_ & new_n_n13_;
  assign new_n_n1076_ = new_n_n16_ & new_nq3_;
  assign new_ny6_ = new_n_n1013_ | new_n_n1011_ | new_n_n1010_ | new_n_n1012_ | new_n_n1014_ | new_n_n1009_ | new_n_n1008_ | new_n_n1007_ | new_n_n1006_;
  assign new_n_n1005_ = new_na17_ & new_nq1_ & new_n_n44_;
  assign new_n_n758_ = new_no0_ & new_n_n189_ & new_n_n188_;
  assign new_n_n722_ = new_nq_ & new_no0_ & new_n_n408_;
  assign new_nj19_ = new_n_n237_ & new_nl4_;
  assign new_nv19_ = new_n_n713_ | new_n_n238_;
  assign new_n_n709_ = new_n_n243_ & new_n_n378_ & new_n_n254_;
  assign new_n_n667_ = new_nk0_ & new_n_n430_ & new_nn_;
  assign new_nc23_ = new_nq2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n604_ = new_n_n330_ & new_ni6_ & new_n_n311_;
  assign new_n_n54_ = ~new_nm18_;
  assign new_n_n43_ = ~new_nl17_;
  assign new_n_n32_ = ~new_nx15_;
  assign new_ng6_ = ~new_nt34_;
  assign new_n_n20_ = ~new_ni34_;
  assign new_n_n14_ = ~new_nv33_;
  assign new_n_n1083_ = new_n_n431_ & new_n_n430_ & new_n_n13_;
  assign new_nz4_ = new_n_n1076_ | new_n_n1075_ | new_n_n1074_;
  assign new_n_n1014_ = new_na17_ & new_np1_ & new_n_n42_;
  assign new_nz6_ = new_n_n1004_ | new_n_n1002_ | new_n_n1001_ | new_n_n1003_ | new_n_n1005_ | new_n_n1000_ | new_n_n999_ | new_n_n998_ | new_n_n997_;
  assign new_nj15_ = new_nc1_ | new_nq0_ | new_n_n411_;
  assign new_nz18_ = new_n_n233_ & new_nl4_;
  assign new_n_n718_ = new_ns_ & new_no0_ & new_n_n408_;
  assign new_n_n713_ = new_n_n239_ & new_n_n378_ & new_n_n254_;
  assign new_nf20_ = new_n_n709_ | new_n_n242_;
  assign new_nu22_ = new_nq2_ | new_n_n365_;
  assign new_nb23_ = new_nr2_ | new_n_n365_;
  assign new_nw16_ = new_n_n387_ & new_nl4_;
  assign new_n_n53_ = ~new_nk18_;
  assign new_n_n44_ = ~new_nn17_;
  assign new_n_n31_ = ~new_ng16_;
  assign new_n_n22_ = ~new_nv34_;
  assign new_nr5_ = ~new_nf34_;
  assign new_n_n15_ = ~new_nw33_;
  assign new_nw4_ = new_n_n1085_ | new_n_n1084_ | new_n_n1083_;
  assign new_n_n1077_ = new_n_n431_ & new_n_n430_ & new_n_n15_;
  assign new_nx15_ = new_n_n378_ | new_ne1_ | new_nn0_;
  assign new_nb19_ = new_n_n721_ | new_n_n230_;
  assign new_n_n717_ = new_n_n235_ & new_n_n378_ & new_n_n254_;
  assign new_n_n714_ = new_nu_ & new_no0_ & new_n_n408_;
  assign new_nd20_ = new_n_n245_ & new_nl4_;
  assign new_n_n679_ = new_nd_ & new_n_n431_;
  assign new_n_n672_ = new_nk0_ & new_n_n430_ & new_nm_;
  assign new_n_n612_ = new_n_n302_ & new_n_n304_ & new_n_n303_;
  assign new_n_n74_ = ~new_nk20_;
  assign new_n_n63_ = ~new_nj19_;
  assign new_n_n30_ = ~new_nb16_;
  assign new_ne6_ = ~new_nr34_;
  assign new_nx5_ = ~new_nk34_;
  assign new_n_n16_ = ~new_nx33_;
  assign new_n_n1085_ = new_n_n13_ & new_nn3_;
  assign new_n_n1078_ = new_nk0_ & new_nl0_ & new_n_n15_;
  assign new_n_n747_ = new_n_n204_ & new_n_n205_;
  assign new_n_n721_ = new_n_n231_ & new_n_n378_ & new_n_n254_;
  assign new_nl19_ = new_n_n717_ | new_n_n234_;
  assign new_nt19_ = new_n_n241_ & new_nl4_;
  assign new_n_n710_ = new_nw_ & new_no0_ & new_n_n408_;
  assign new_n_n678_ = new_nd_ & new_nl0_;
  assign new_n_n673_ = new_ne_ & new_nl0_;
  assign new_n_n619_ = new_n_n298_ & new_na17_ & new_n_n299_;
  assign new_n_n73_ = ~new_ni20_;
  assign new_n_n64_ = ~new_nl19_;
  assign new_n_n29_ = ~new_nc16_;
  assign new_nf6_ = ~new_ns34_;
  assign new_n_n21_ = ~new_nh34_;
  assign new_n_n17_ = ~new_ny33_;
  assign new_n_n1079_ = new_n_n15_ & new_np3_;
  assign new_ns16_ = new_nn0_ | new_n_n378_;
  assign new_n_n706_ = new_ny_ & new_no0_ & new_n_n408_;
  assign new_nx20_ = new_n_n255_ & new_nl4_;
  assign new_nh21_ = new_n_n256_ | new_n_n696_ | new_n_n695_;
  assign new_n_n691_ = new_n_n428_ & new_n_n350_ & new_n_n260_;
  assign new_n_n690_ = new_n_n387_ & new_n_n261_ & new_n_n279_;
  assign new_n_n684_ = new_nc_ & new_n_n431_;
  assign new_n_n626_ = new_n_n296_ & new_n_n301_;
  assign new_n_n75_ = ~new_nn20_;
  assign new_n_n72_ = ~new_nf20_;
  assign new_n_n61_ = ~new_ne19_;
  assign new_n_n50_ = ~new_nc18_;
  assign new_n_n39_ = ~new_nb17_;
  assign new_nz5_ = ~new_nm34_;
  assign new_n_n18_ = ~new_nz33_;
  assign new_n_n1086_ = new_n_n431_ & new_n_n430_ & new_n_n12_;
  assign new_n_n741_ = new_n_n211_ & new_n_n378_ & new_n_n254_;
  assign new_nn20_ = new_n_n249_ & new_nl4_;
  assign new_n_n702_ = new_na0_ & new_no0_ & new_n_n408_;
  assign new_n_n696_ = new_n_n428_ & new_n_n350_ & new_n_n257_;
  assign new_nq21_ = new_n_n259_ | new_n_n691_ | new_n_n690_;
  assign new_nr21_ = new_n_n689_ | new_n_n688_ | new_n_n687_;
  assign new_ny21_ = new_n_n684_ | new_n_n683_ | new_n_n682_;
  assign new_ng24_ = new_n_n629_ | new_n_n631_ | new_n_n630_ | new_n_n632_;
  assign new_n_n76_ = ~new_np20_;
  assign new_n_n71_ = ~new_nd20_;
  assign new_n_n62_ = ~new_ng19_;
  assign new_n_n49_ = ~new_na18_;
  assign new_n_n40_ = ~new_nd17_;
  assign new_ny5_ = ~new_nl34_;
  assign new_n_n19_ = ~new_na34_;
  assign new_n_n737_ = new_n_n215_ & new_n_n378_ & new_n_n254_;
  assign new_np20_ = new_n_n705_ | new_n_n246_;
  assign new_n_n701_ = new_n_n251_ & new_n_n378_ & new_n_n254_;
  assign new_n_n698_ = new_nc0_ & new_no0_ & new_n_n408_;
  assign new_nl21_ = new_nk2_ | new_n_n656_ | new_n_n655_;
  assign new_n_n77_ = ~new_ns20_;
  assign new_n_n70_ = ~new_na20_;
  assign new_n_n59_ = ~new_nz18_;
  assign new_n_n52_ = ~new_nh18_;
  assign new_n_n41_ = ~new_ng17_;
  assign new_n_n34_ = ~new_nj16_;
  assign new_n_n23_ = ~new_nk15_;
  assign new_n_n733_ = new_n_n219_ & new_n_n378_ & new_n_n254_;
  assign new_n_n705_ = new_n_n247_ & new_n_n378_ & new_n_n254_;
  assign new_nz20_ = new_n_n701_ | new_n_n250_;
  assign new_n_n697_ = new_n_n378_ & new_no0_ & new_n_n408_;
  assign new_nk21_ = new_nt15_ & new_n_n432_ & new_n_n428_;
  assign new_n_n78_ = ~new_nu20_;
  assign new_n_n69_ = ~new_ny19_;
  assign new_n_n60_ = ~new_nb19_;
  assign new_n_n51_ = ~new_nf18_;
  assign new_n_n42_ = ~new_ni17_;
  assign new_n_n33_ = ~new_nf16_;
  assign new_n_n24_ = ~new_nj15_;
endmodule


