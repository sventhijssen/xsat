// Benchmark "top" written by ABC on Fri Mar 31 12:07:32 2023

module top ( 
    i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_, i_10_,
    i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_,
    i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_, i_24_,
    i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_, i_32_,
    i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_, i_19_,
    i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_, i_38_,
    i_29_, i_51_, i_44_, i_37_,
    o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_  );
  input  i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_,
    i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_,
    i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_,
    i_24_, i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_,
    i_32_, i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_,
    i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_,
    i_38_, i_29_, i_51_, i_44_, i_37_;
  output o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_;
  wire new_ni_63__, new_ni_50__, new_ni_64__, new_ni_61__, new_ni_62__,
    new_ni_40__, new_ni_30__, new_ni_20__, new_ni_9__, new_ni_10__,
    new_ni_7__, new_ni_8__, new_ni_5__, new_ni_6__, new_ni_27__,
    new_ni_14__, new_ni_3__, new_ni_39__, new_ni_28__, new_ni_13__,
    new_ni_4__, new_ni_25__, new_ni_12__, new_ni_1__, new_ni_26__,
    new_ni_11__, new_ni_2__, new_ni_49__, new_ni_23__, new_ni_18__,
    new_ni_24__, new_ni_17__, new_ni_0__, new_ni_21__, new_ni_16__,
    new_ni_59__, new_ni_22__, new_ni_15__, new_ni_58__, new_ni_45__,
    new_ni_32__, new_ni_57__, new_ni_46__, new_ni_31__, new_ni_56__,
    new_ni_47__, new_ni_34__, new_ni_55__, new_ni_48__, new_ni_33__,
    new_ni_19__, new_ni_54__, new_ni_41__, new_ni_36__, new_ni_60__,
    new_ni_53__, new_ni_42__, new_ni_35__, new_ni_52__, new_ni_43__,
    new_ni_38__, new_ni_29__, new_ni_51__, new_ni_44__, new_ni_37__,
    new_no_4__, new_n_n449_, new_n_n438_, new_n_n427_, new_n_n416_,
    new_n_n405_, new_n_n394_, new_no_63__, new_n_n375_, new_n_n366_,
    new_n_n356_, new_no_57__, new_n_n325_, new_n_n315_, new_n_n306_,
    new_no_53__, new_n_n285_, new_n_n275_, new_n_n266_, new_n_n256_,
    new_n_n227_, new_n_n217_, new_n_n208_, new_n_n198_, new_n_n189_,
    new_n_n179_, new_no_36__, new_n_n134_, new_n_n124_, new_n_n114_,
    new_n_n105_, new_n_n95_, new_n_n86_, new_n_n448_, new_n_n439_,
    new_n_n437_, new_n_n415_, new_n_n406_, new_n_n393_, new_n_n385_,
    new_n_n374_, new_no_60__, new_n_n355_, new_n_n347_, new_n_n324_,
    new_n_n316_, new_n_n305_, new_n_n296_, new_n_n284_, new_n_n276_,
    new_n_n265_, new_n_n257_, new_n_n236_, new_n_n216_, new_n_n209_,
    new_n_n197_, new_n_n190_, new_n_n178_, new_n_n170_, new_n_n133_,
    new_n_n125_, new_n_n113_, new_n_n106_, new_n_n94_, new_no_21__,
    new_n_n458_, new_n_n451_, new_n_n440_, new_n_n414_, new_n_n403_,
    new_n_n396_, new_n_n386_, new_no_61__, new_n_n364_, new_n_n358_,
    new_n_n348_, new_n_n323_, new_n_n313_, new_n_n307_, new_n_n297_,
    new_n_n283_, new_n_n274_, new_n_n268_, new_n_n258_, new_n_n235_,
    new_n_n225_, new_no_42__, new_no_40__, new_n_n187_, new_n_n181_,
    new_n_n171_, new_no_31__, new_n_n141_, new_n_n112_, new_n_n103_,
    new_n_n97_, new_n_n87_, new_no_11__, new_n_n450_, new_n_n441_,
    new_n_n413_, new_n_n404_, new_n_n395_, new_n_n387_, new_n_n373_,
    new_n_n365_, new_n_n357_, new_n_n349_, new_n_n322_, new_n_n314_,
    new_no_54__, new_n_n298_, new_n_n282_, new_no_51__, new_n_n267_,
    new_n_n259_, new_n_n234_, new_n_n226_, new_n_n218_, new_n_n196_,
    new_n_n188_, new_n_n180_, new_n_n172_, new_n_n150_, new_n_n142_,
    new_no_25__, new_n_n104_, new_n_n96_, new_n_n88_, new_n_n434_,
    new_n_n423_, new_no_64__, new_n_n372_, new_n_n343_, new_n_n332_,
    new_n_n281_, new_n_n272_, new_n_n253_, new_n_n243_, new_n_n195_,
    new_n_n186_, new_n_n175_, new_n_n166_, new_no_33__, new_n_n111_,
    new_n_n101_, new_n_n91_, new_no_20__, new_n_n8_, new_n_n433_,
    new_n_n424_, new_n_n397_, new_n_n363_, new_n_n342_, new_n_n333_,
    new_n_n280_, new_n_n273_, new_n_n252_, new_n_n244_, new_n_n194_,
    new_no_38__, new_n_n167_, new_n_n165_, new_n_n158_, new_n_n110_,
    new_n_n102_, new_no_22__, new_n_n83_, new_n_n436_, new_n_n425_,
    new_n_n407_, new_no_58__, new_n_n345_, new_n_n334_, new_n_n264_,
    new_n_n254_, new_n_n245_, new_n_n193_, new_n_n177_, new_n_n168_,
    new_n_n109_, new_n_n99_, new_n_n93_, new_n_n84_, new_n_n435_,
    new_n_n426_, new_n_n417_, new_n_n346_, new_n_n344_, new_n_n335_,
    new_n_n263_, new_n_n255_, new_no_48__, new_n_n185_, new_n_n176_,
    new_n_n169_, new_n_n108_, new_n_n100_, new_n_n92_, new_n_n85_,
    new_n_n457_, new_n_n446_, new_n_n430_, new_n_n419_, new_n_n408_,
    new_n_n354_, new_n_n339_, new_n_n328_, new_n_n318_, new_n_n308_,
    new_n_n249_, new_no_46__, new_n_n230_, new_no_44__, new_n_n210_,
    new_n_n162_, new_n_n155_, new_n_n145_, new_n_n137_, new_n_n127_,
    new_no_26__, new_n_n4_, new_n_n456_, new_n_n447_, new_n_n429_,
    new_n_n420_, new_n_n398_, new_no_59__, new_n_n338_, new_n_n329_,
    new_n_n317_, new_n_n309_, new_n_n248_, new_n_n240_, new_n_n229_,
    new_n_n220_, new_n_n202_, new_no_35__, new_n_n156_, new_n_n144_,
    new_no_28__, new_n_n126_, new_n_n117_, new_n_n5_, new_n_n432_,
    new_n_n421_, new_n_n388_, new_n_n371_, new_n_n341_, new_n_n330_,
    new_n_n300_, new_n_n290_, new_n_n251_, new_n_n241_, new_n_n228_,
    new_n_n212_, new_n_n203_, new_n_n164_, new_no_32__, new_n_n143_,
    new_n_n135_, new_no_27__, new_n_n118_, new_n_n6_, new_n_n431_,
    new_n_n422_, new_no_62__, new_n_n380_, new_n_n340_, new_n_n331_,
    new_n_n299_, new_n_n291_, new_n_n250_, new_n_n242_, new_n_n219_,
    new_n_n211_, new_no_41__, new_n_n163_, new_n_n157_, new_no_30__,
    new_n_n136_, new_n_n128_, new_n_n119_, new_n_n7_, new_n_n453_,
    new_n_n442_, new_n_n412_, new_n_n401_, new_n_n390_, new_n_n381_,
    new_n_n379_, new_n_n369_, new_n_n360_, new_n_n350_, new_no_56__,
    new_n_n311_, new_n_n302_, new_n_n292_, new_n_n289_, new_n_n279_,
    new_n_n269_, new_no_49__, new_no_47__, new_n_n233_, new_n_n223_,
    new_no_43__, new_n_n204_, new_n_n192_, new_n_n183_, new_n_n173_,
    new_n_n160_, new_n_n151_, new_n_n149_, new_n_n140_, new_n_n130_,
    new_n_n120_, new_n_n98_, new_n_n89_, new_n_n0_, new_n_n452_,
    new_n_n443_, new_n_n411_, new_n_n402_, new_n_n389_, new_n_n382_,
    new_n_n378_, new_n_n370_, new_n_n359_, new_n_n351_, new_n_n321_,
    new_n_n312_, new_n_n301_, new_n_n293_, new_n_n288_, new_no_52__,
    new_no_50__, new_n_n260_, new_n_n237_, new_n_n232_, new_n_n224_,
    new_n_n213_, new_n_n205_, new_n_n201_, new_n_n182_, new_no_37__,
    new_n_n159_, new_n_n152_, new_n_n148_, new_no_29__, new_n_n129_,
    new_n_n121_, new_no_23__, new_n_n90_, new_n_n1_, new_n_n455_,
    new_n_n444_, new_n_n428_, new_n_n410_, new_n_n399_, new_n_n392_,
    new_n_n383_, new_n_n377_, new_n_n367_, new_n_n362_, new_n_n352_,
    new_n_n337_, new_n_n326_, new_n_n320_, new_n_n310_, new_n_n304_,
    new_n_n294_, new_n_n287_, new_n_n277_, new_n_n271_, new_n_n261_,
    new_n_n247_, new_n_n238_, new_no_45__, new_n_n221_, new_n_n215_,
    new_n_n206_, new_n_n200_, new_no_39__, new_n_n174_, new_n_n161_,
    new_n_n153_, new_n_n147_, new_n_n138_, new_n_n132_, new_n_n122_,
    new_n_n116_, new_n_n107_, new_n_n2_, new_n_n454_, new_n_n445_,
    new_n_n418_, new_n_n409_, new_n_n400_, new_n_n391_, new_n_n384_,
    new_n_n376_, new_n_n368_, new_n_n361_, new_n_n353_, new_n_n336_,
    new_n_n327_, new_n_n319_, new_no_55__, new_n_n303_, new_n_n295_,
    new_n_n286_, new_n_n278_, new_n_n270_, new_n_n262_, new_n_n246_,
    new_n_n239_, new_n_n231_, new_n_n222_, new_n_n214_, new_n_n207_,
    new_n_n199_, new_n_n191_, new_n_n184_, new_no_34__, new_n_n154_,
    new_n_n146_, new_n_n139_, new_n_n131_, new_n_n123_, new_n_n115_,
    new_no_24__, new_n_n3_, new_n_n78_, new_n_n69_, new_n_n61_, new_n_n53_,
    new_n_n43_, new_no_19__, new_n_n68_, new_n_n62_, new_n_n52_,
    new_n_n44_, new_n_n79_, new_no_16__, new_no_13__, new_n_n54_,
    new_no_9__, new_n_n80_, new_n_n67_, new_n_n60_, new_no_10__,
    new_n_n45_, new_no_0__, new_n_n81_, new_n_n37_, new_n_n28_, new_n_n18_,
    new_n_n9_, new_n_n82_, new_n_n36_, new_n_n29_, new_n_n17_, new_no_1__,
    new_no_7__, new_n_n26_, new_n_n20_, new_n_n10_, new_n_n35_, new_n_n27_,
    new_n_n19_, new_n_n11_, new_n_n59_, new_n_n50_, new_n_n40_, new_n_n32_,
    new_n_n22_, new_n_n12_, new_n_n58_, new_n_n51_, new_n_n39_, new_n_n33_,
    new_n_n21_, new_n_n13_, new_n_n74_, new_no_15__, new_n_n38_,
    new_n_n30_, new_n_n24_, new_n_n14_, new_n_n73_, new_n_n66_, new_no_8__,
    new_n_n31_, new_n_n23_, new_n_n15_, new_no_18__, new_n_n72_,
    new_no_14__, new_n_n55_, new_n_n46_, new_no_3__, new_no_2__,
    new_n_n75_, new_n_n71_, new_n_n65_, new_no_12__, new_n_n47_,
    new_n_n25_, new_n_n16_, new_n_n76_, new_no_17__, new_n_n63_,
    new_n_n57_, new_n_n48_, new_n_n42_, new_no_6__, new_n_n77_, new_n_n70_,
    new_n_n64_, new_n_n56_, new_n_n49_, new_n_n41_, new_n_n34_;
  assign o_1_ = new_no_1__;
  assign new_ni_63__ = i_63_;
  assign new_ni_50__ = i_50_;
  assign o_19_ = new_no_19__;
  assign o_2_ = new_no_2__;
  assign new_ni_64__ = i_64_;
  assign new_ni_61__ = i_61_;
  assign o_0_ = new_no_0__;
  assign new_ni_62__ = i_62_;
  assign new_ni_40__ = i_40_;
  assign o_29_ = new_no_29__;
  assign new_ni_30__ = i_30_;
  assign o_60_ = new_no_60__;
  assign o_39_ = new_no_39__;
  assign o_38_ = new_no_38__;
  assign o_25_ = new_no_25__;
  assign o_12_ = new_no_12__;
  assign o_37_ = new_no_37__;
  assign o_26_ = new_no_26__;
  assign o_11_ = new_no_11__;
  assign new_ni_20__ = i_20_;
  assign o_50_ = new_no_50__;
  assign o_36_ = new_no_36__;
  assign o_27_ = new_no_27__;
  assign o_14_ = new_no_14__;
  assign new_ni_9__ = i_9_;
  assign o_35_ = new_no_35__;
  assign o_28_ = new_no_28__;
  assign o_13_ = new_no_13__;
  assign o_34_ = new_no_34__;
  assign o_21_ = new_no_21__;
  assign o_16_ = new_no_16__;
  assign new_ni_10__ = i_10_;
  assign new_ni_7__ = i_7_;
  assign o_40_ = new_no_40__;
  assign o_33_ = new_no_33__;
  assign o_22_ = new_no_22__;
  assign o_15_ = new_no_15__;
  assign new_ni_8__ = i_8_;
  assign o_32_ = new_no_32__;
  assign o_23_ = new_no_23__;
  assign o_18_ = new_no_18__;
  assign new_ni_5__ = i_5_;
  assign o_31_ = new_no_31__;
  assign o_24_ = new_no_24__;
  assign o_17_ = new_no_17__;
  assign new_ni_6__ = i_6_;
  assign o_56_ = new_no_56__;
  assign o_43_ = new_no_43__;
  assign o_30_ = new_no_30__;
  assign new_ni_27__ = i_27_;
  assign new_ni_14__ = i_14_;
  assign new_ni_3__ = i_3_;
  assign o_55_ = new_no_55__;
  assign o_44_ = new_no_44__;
  assign new_ni_39__ = i_39_;
  assign new_ni_28__ = i_28_;
  assign new_ni_13__ = i_13_;
  assign new_ni_4__ = i_4_;
  assign o_58_ = new_no_58__;
  assign o_41_ = new_no_41__;
  assign new_ni_25__ = i_25_;
  assign new_ni_12__ = i_12_;
  assign new_ni_1__ = i_1_;
  assign o_57_ = new_no_57__;
  assign o_42_ = new_no_42__;
  assign o_20_ = new_no_20__;
  assign new_ni_26__ = i_26_;
  assign new_ni_11__ = i_11_;
  assign new_ni_2__ = i_2_;
  assign o_52_ = new_no_52__;
  assign o_47_ = new_no_47__;
  assign new_ni_49__ = i_49_;
  assign new_ni_23__ = i_23_;
  assign new_ni_18__ = i_18_;
  assign o_51_ = new_no_51__;
  assign o_48_ = new_no_48__;
  assign new_ni_24__ = i_24_;
  assign new_ni_17__ = i_17_;
  assign new_ni_0__ = i_0_;
  assign o_54_ = new_no_54__;
  assign o_45_ = new_no_45__;
  assign o_10_ = new_no_10__;
  assign new_ni_21__ = i_21_;
  assign new_ni_16__ = i_16_;
  assign o_53_ = new_no_53__;
  assign o_46_ = new_no_46__;
  assign new_ni_59__ = i_59_;
  assign new_ni_22__ = i_22_;
  assign new_ni_15__ = i_15_;
  assign o_61_ = new_no_61__;
  assign o_9_ = new_no_9__;
  assign new_ni_58__ = i_58_;
  assign new_ni_45__ = i_45_;
  assign new_ni_32__ = i_32_;
  assign o_62_ = new_no_62__;
  assign new_ni_57__ = i_57_;
  assign new_ni_46__ = i_46_;
  assign new_ni_31__ = i_31_;
  assign o_63_ = new_no_63__;
  assign o_49_ = new_no_49__;
  assign o_7_ = new_no_7__;
  assign new_ni_56__ = i_56_;
  assign new_ni_47__ = i_47_;
  assign new_ni_34__ = i_34_;
  assign o_64_ = new_no_64__;
  assign o_8_ = new_no_8__;
  assign new_ni_55__ = i_55_;
  assign new_ni_48__ = i_48_;
  assign new_ni_33__ = i_33_;
  assign new_ni_19__ = i_19_;
  assign o_5_ = new_ni_29__;
  assign new_ni_54__ = i_54_;
  assign new_ni_41__ = i_41_;
  assign new_ni_36__ = i_36_;
  assign o_59_ = new_no_59__;
  assign o_6_ = new_no_6__;
  assign new_ni_60__ = i_60_;
  assign new_ni_53__ = i_53_;
  assign new_ni_42__ = i_42_;
  assign new_ni_35__ = i_35_;
  assign o_3_ = new_no_3__;
  assign new_ni_52__ = i_52_;
  assign new_ni_43__ = i_43_;
  assign new_ni_38__ = i_38_;
  assign new_ni_29__ = i_29_;
  assign o_4_ = new_no_4__;
  assign new_ni_51__ = i_51_;
  assign new_ni_44__ = i_44_;
  assign new_ni_37__ = i_37_;
  assign new_no_4__ = new_ni_29__ & new_ni_15__;
  assign new_n_n449_ = ~new_ni_40__;
  assign new_n_n438_ = ~new_ni_6__;
  assign new_n_n427_ = ~new_ni_9__;
  assign new_n_n416_ = ~new_ni_42__;
  assign new_n_n405_ = ~new_ni_61__;
  assign new_n_n394_ = new_n_n455_ & new_n_n454_ & new_n_n453_;
  assign new_no_63__ = new_n_n385_ & new_n_n382_;
  assign new_n_n375_ = new_n_n380_ & new_n_n58_ & new_n_n379_;
  assign new_n_n366_ = new_n_n458_ & new_n_n456_ & new_n_n455_;
  assign new_n_n356_ = new_n_n360_ & new_n_n387_ & new_n_n392_;
  assign new_no_57__ = new_n_n434_ & new_n_n347_;
  assign new_n_n325_ = new_n_n334_ & new_n_n333_ & new_n_n332_;
  assign new_n_n315_ = new_n_n321_ & new_n_n320_ & new_n_n372_;
  assign new_n_n306_ = new_n_n456_ & new_n_n455_ & new_n_n424_;
  assign new_no_53__ = new_n_n296_ & new_n_n297_;
  assign new_n_n285_ = new_n_n403_ & new_n_n404_;
  assign new_n_n275_ = new_n_n271_ & new_n_n276_ & new_n_n206_;
  assign new_n_n266_ = new_n_n416_ & new_n_n448_ & new_n_n447_;
  assign new_n_n256_ = new_n_n278_ & new_n_n277_ & new_n_n434_;
  assign new_n_n227_ = new_n_n443_ & new_n_n421_ & new_n_n420_;
  assign new_n_n217_ = new_n_n343_ & new_n_n306_ & new_n_n319_;
  assign new_n_n208_ = new_n_n209_ & new_n_n267_ & new_n_n338_;
  assign new_n_n198_ = new_n_n263_ & new_n_n236_ & new_n_n201_;
  assign new_n_n189_ = new_n_n293_ & new_n_n292_ & new_n_n238_;
  assign new_n_n179_ = new_n_n305_ & new_n_n183_ & new_n_n182_;
  assign new_no_36__ = new_n_n171_ & new_n_n170_;
  assign new_n_n134_ = new_n_n227_ & new_n_n155_ & new_n_n392_;
  assign new_n_n124_ = new_n_n434_ & new_n_n404_ & new_n_n403_;
  assign new_n_n114_ = new_n_n446_ & new_n_n445_ & new_n_n444_;
  assign new_n_n105_ = new_n_n417_ & new_n_n451_ & new_n_n450_;
  assign new_n_n95_ = new_n_n360_ & new_n_n387_ & new_n_n339_;
  assign new_n_n86_ = new_n_n446_ & new_ni_51__ & new_n_n442_;
  assign new_n_n448_ = ~new_ni_43__;
  assign new_n_n439_ = ~new_ni_3__;
  assign new_n_n437_ = ~new_ni_7__;
  assign new_n_n415_ = ~new_ni_45__;
  assign new_n_n406_ = ~new_ni_59__;
  assign new_n_n393_ = new_n_n452_ & new_ni_29__ & new_ni_30__;
  assign new_n_n385_ = new_n_n392_ & new_n_n391_ & new_n_n386_;
  assign new_n_n374_ = new_n_n378_ & new_n_n377_ & new_n_n376_;
  assign new_no_60__ = new_n_n367_ & new_n_n76_ & new_n_n368_;
  assign new_n_n355_ = new_n_n359_ & new_n_n376_ & new_n_n358_;
  assign new_n_n347_ = new_n_n350_ & new_n_n349_ & new_n_n348_;
  assign new_n_n324_ = new_n_n403_ & new_n_n331_;
  assign new_n_n316_ = new_n_n441_ & new_n_n446_ & new_n_n412_;
  assign new_n_n305_ = new_ni_29__ & new_n_n443_ & new_n_n421_;
  assign new_n_n296_ = new_n_n271_ & new_n_n81_ & new_n_n298_;
  assign new_n_n284_ = new_n_n343_ & new_n_n295_ & new_n_n294_;
  assign new_n_n276_ = new_n_n279_ & new_n_n300_ & new_n_n278_;
  assign new_n_n265_ = new_ni_53__ & new_n_n409_ & new_n_n408_;
  assign new_n_n257_ = new_n_n303_ & new_n_n369_ & new_n_n300_;
  assign new_n_n236_ = new_n_n306_ & new_n_n319_ & new_n_n318_;
  assign new_n_n216_ = new_n_n289_ & new_n_n288_ & new_n_n332_;
  assign new_n_n209_ = new_ni_29__ & new_n_n443_ & new_ni_33__;
  assign new_n_n197_ = new_n_n199_ & new_n_n200_;
  assign new_n_n190_ = new_n_n442_ & new_n_n445_ & new_ni_59__;
  assign new_n_n178_ = new_n_n338_ & new_n_n337_ & new_n_n336_;
  assign new_n_n170_ = new_n_n315_ & new_n_n172_ & new_n_n313_;
  assign new_n_n133_ = new_n_n303_ & new_n_n302_ & new_n_n301_;
  assign new_n_n125_ = new_n_n442_ & new_n_n407_ & new_n_n445_;
  assign new_n_n113_ = new_n_n366_ & new_n_n116_ & new_n_n115_;
  assign new_n_n106_ = new_n_n422_ & new_n_n433_ & new_n_n454_;
  assign new_n_n94_ = new_n_n97_ & new_n_n338_ & new_n_n337_;
  assign new_no_21__ = new_n_n308_ & new_n_n87_;
  assign new_n_n458_ = ~new_ni_10__;
  assign new_n_n451_ = ~new_ni_37__;
  assign new_n_n440_ = ~new_ni_8__;
  assign new_n_n414_ = ~new_ni_48__;
  assign new_n_n403_ = ~new_ni_64__;
  assign new_n_n396_ = ~new_ni_44__;
  assign new_n_n386_ = new_ni_56__ & new_n_n445_ & new_n_n444_;
  assign new_no_61__ = new_n_n375_ & new_n_n374_ & new_n_n390_;
  assign new_n_n364_ = new_ni_40__ & new_n_n448_ & new_n_n446_;
  assign new_n_n358_ = new_n_n445_ & new_n_n444_ & new_n_n434_;
  assign new_n_n348_ = new_n_n168_ & new_n_n369_ & new_n_n368_;
  assign new_n_n323_ = new_n_n330_ & new_n_n329_ & new_n_n328_;
  assign new_n_n313_ = new_n_n392_ & new_n_n359_ & new_n_n316_;
  assign new_n_n307_ = new_n_n308_ & new_n_n309_;
  assign new_n_n297_ = new_n_n330_ & new_n_n217_ & new_n_n272_;
  assign new_n_n283_ = new_n_n293_ & new_n_n292_ & new_n_n291_;
  assign new_n_n274_ = new_n_n408_ & new_n_n442_ & new_ni_57__;
  assign new_n_n268_ = new_n_n432_ & new_n_n439_ & new_n_n429_;
  assign new_n_n258_ = new_n_n259_ & new_n_n304_ & new_n_n392_;
  assign new_n_n235_ = new_n_n239_ & new_n_n293_ & new_n_n292_;
  assign new_n_n225_ = new_n_n395_ & new_n_n228_ & new_n_n352_;
  assign new_no_42__ = new_n_n210_ & new_n_n297_;
  assign new_no_40__ = new_n_n197_ & new_n_n198_;
  assign new_n_n187_ = new_n_n251_ & new_n_n194_ & new_n_n189_;
  assign new_n_n181_ = new_n_n343_ & new_n_n186_ & new_n_n185_;
  assign new_n_n171_ = new_n_n173_ & new_n_n278_;
  assign new_no_31__ = new_n_n152_ & new_n_n151_ & new_n_n403_;
  assign new_n_n141_ = new_ni_60__ & new_n_n110_;
  assign new_n_n112_ = new_n_n114_ & new_n_n377_;
  assign new_n_n103_ = new_n_n106_ & new_n_n318_ & new_n_n305_;
  assign new_n_n97_ = new_n_n418_ & new_ni_36__ & new_n_n451_;
  assign new_n_n87_ = new_n_n89_ & new_n_n85_ & new_n_n88_;
  assign new_no_11__ = new_n_n455_ & new_ni_29__ & new_ni_37__;
  assign new_n_n450_ = ~new_ni_39__;
  assign new_n_n441_ = ~new_ni_47__;
  assign new_n_n413_ = ~new_ni_49__;
  assign new_n_n404_ = ~new_ni_63__;
  assign new_n_n395_ = new_n_n458_ & new_n_n457_ & new_n_n456_;
  assign new_n_n387_ = new_n_n452_ & new_ni_29__ & new_n_n443_;
  assign new_n_n373_ = new_ni_7__ & new_n_n440_ & new_n_n458_;
  assign new_n_n365_ = new_n_n452_ & new_ni_29__ & new_n_n451_;
  assign new_n_n357_ = new_n_n354_ & new_n_n362_ & new_n_n361_;
  assign new_n_n349_ = new_n_n352_ & new_n_n351_ & new_n_n378_;
  assign new_n_n322_ = new_n_n327_ & new_n_n326_ & new_n_n325_;
  assign new_n_n314_ = new_n_n319_ & new_n_n318_ & new_n_n317_;
  assign new_no_54__ = new_n_n307_ & new_n_n170_;
  assign new_n_n298_ = new_n_n332_ & new_n_n299_ & new_n_n403_;
  assign new_n_n282_ = new_n_n290_ & new_n_n289_ & new_n_n288_;
  assign new_no_51__ = new_n_n275_ & new_n_n297_;
  assign new_n_n267_ = new_n_n419_ & new_n_n418_ & new_n_n451_;
  assign new_n_n259_ = new_ni_29__ & new_n_n443_ & new_ni_31__;
  assign new_n_n234_ = new_n_n238_ & new_n_n237_ & new_n_n264_;
  assign new_n_n226_ = new_n_n231_ & new_n_n230_ & new_n_n229_;
  assign new_n_n218_ = new_n_n219_ & new_n_n345_ & new_n_n344_;
  assign new_n_n196_ = new_n_n455_ & new_n_n423_ & new_n_n433_;
  assign new_n_n188_ = new_n_n237_ & new_n_n190_ & new_n_n286_;
  assign new_n_n180_ = new_n_n184_ & new_n_n106_ & new_n_n318_;
  assign new_n_n172_ = new_n_n319_ & new_n_n318_ & new_n_n310_;
  assign new_n_n150_ = new_n_n424_ & new_n_n423_ & new_n_n422_;
  assign new_n_n142_ = new_n_n366_ & new_n_n365_ & new_n_n370_;
  assign new_no_25__ = new_n_n112_ & new_n_n113_;
  assign new_n_n104_ = new_n_n343_ & new_n_n342_ & new_n_n107_;
  assign new_n_n96_ = new_n_n343_ & new_n_n342_ & new_n_n294_;
  assign new_n_n88_ = new_n_n338_ & new_n_n238_ & new_n_n383_;
  assign new_n_n434_ = ~new_ni_62__;
  assign new_n_n423_ = ~new_ni_18__;
  assign new_no_64__ = new_n_n388_ & new_n_n389_;
  assign new_n_n372_ = new_n_n457_ & new_n_n456_ & new_n_n455_;
  assign new_n_n343_ = new_n_n427_ & new_n_n458_ & new_n_n457_;
  assign new_n_n332_ = new_n_n445_ & new_n_n406_ & new_n_n444_;
  assign new_n_n281_ = new_n_n330_ & new_n_n284_ & new_n_n95_;
  assign new_n_n272_ = new_n_n318_ & new_n_n305_ & new_n_n304_;
  assign new_n_n253_ = new_n_n455_ & new_ni_17__ & new_n_n423_;
  assign new_n_n243_ = new_n_n310_ & new_n_n392_ & new_n_n303_;
  assign new_n_n195_ = new_n_n449_ & new_n_n435_ & new_ni_42__;
  assign new_n_n186_ = new_n_n426_ & new_n_n402_ & new_n_n456_;
  assign new_n_n175_ = new_n_n330_ & new_n_n181_ & new_n_n180_;
  assign new_n_n166_ = new_n_n445_ & new_n_n444_ & new_n_n405_;
  assign new_no_33__ = new_n_n159_ & new_n_n158_;
  assign new_n_n111_ = new_n_n458_ & new_ni_11__ & new_n_n456_;
  assign new_n_n101_ = new_n_n291_ & new_n_n290_ & new_n_n126_;
  assign new_n_n91_ = new_n_n94_ & new_n_n93_ & new_n_n40_;
  assign new_no_20__ = new_n_n358_ & new_n_n83_;
  assign new_n_n8_ = new_n_n440_ & new_n_n427_ & new_n_n458_;
  assign new_n_n433_ = ~new_ni_22__;
  assign new_n_n424_ = ~new_ni_17__;
  assign new_n_n397_ = ~new_ni_38__;
  assign new_n_n363_ = new_n_n366_ & new_n_n365_ & new_n_n364_;
  assign new_n_n342_ = new_n_n426_ & new_n_n456_ & new_n_n455_;
  assign new_n_n333_ = new_n_n408_ & new_n_n442_ & new_n_n407_;
  assign new_n_n280_ = new_n_n283_ & new_n_n282_ & new_n_n47_;
  assign new_n_n273_ = new_n_n434_ & new_n_n405_;
  assign new_n_n252_ = new_n_n443_ & new_n_n418_ & new_n_n451_;
  assign new_n_n244_ = new_n_n268_ & new_n_n344_ & new_n_n245_;
  assign new_n_n194_ = new_n_n196_ & new_n_n360_ & new_n_n387_;
  assign new_no_38__ = new_n_n188_ & new_n_n187_;
  assign new_n_n167_ = new_n_n412_ & new_n_n408_ & new_n_n442_;
  assign new_n_n165_ = new_n_n169_ & new_n_n344_ & new_n_n395_;
  assign new_n_n158_ = new_n_n366_ & new_n_n365_ & new_n_n160_;
  assign new_n_n110_ = new_n_n447_ & new_n_n446_ & new_n_n445_;
  assign new_n_n102_ = new_n_n304_ & new_n_n105_ & new_n_n292_;
  assign new_no_22__ = new_n_n91_ & new_n_n92_;
  assign new_n_n83_ = new_n_n315_ & new_n_n85_ & new_n_n84_;
  assign new_n_n436_ = ~new_ni_26__;
  assign new_n_n425_ = ~new_ni_16__;
  assign new_n_n407_ = ~new_ni_57__;
  assign new_no_58__ = new_n_n357_ & new_n_n356_ & new_n_n355_;
  assign new_n_n345_ = new_n_n439_ & new_n_n429_ & new_n_n428_;
  assign new_n_n334_ = new_n_n411_ & new_n_n410_ & new_n_n409_;
  assign new_n_n264_ = new_n_n442_ & new_n_n445_ & new_n_n406_;
  assign new_n_n254_ = new_n_n256_ & new_n_n257_;
  assign new_n_n245_ = new_ni_9__ & new_n_n458_ & new_n_n457_;
  assign new_n_n193_ = new_n_n293_ & new_n_n195_ & new_n_n238_;
  assign new_n_n177_ = new_n_n335_ & new_n_n334_ & new_n_n333_;
  assign new_n_n168_ = new_n_n449_ & new_n_n435_ & new_n_n448_;
  assign new_n_n109_ = new_n_n111_ & new_n_n394_ & new_n_n365_;
  assign new_n_n99_ = new_n_n330_ & new_n_n104_ & new_n_n103_;
  assign new_n_n93_ = new_n_n336_ & new_n_n335_ & new_n_n212_;
  assign new_n_n84_ = new_n_n338_ & new_n_n238_ & new_n_n86_;
  assign new_n_n435_ = ~new_ni_41__;
  assign new_n_n426_ = ~new_ni_12__;
  assign new_n_n417_ = ~new_ni_36__;
  assign new_n_n346_ = new_n_n432_ & new_n_n431_ & new_n_n430_;
  assign new_n_n344_ = new_n_n438_ & new_n_n437_ & new_n_n440_;
  assign new_n_n335_ = new_n_n413_ & new_n_n446_ & new_n_n412_;
  assign new_n_n263_ = new_n_n268_ & new_n_n344_ & new_n_n343_;
  assign new_n_n255_ = new_n_n263_ & new_n_n236_ & new_n_n258_;
  assign new_no_48__ = new_n_n254_ & new_n_n255_;
  assign new_n_n185_ = new_n_n455_ & new_n_n425_ & new_n_n424_;
  assign new_n_n176_ = new_n_n332_ & new_n_n331_ & new_n_n403_;
  assign new_n_n169_ = new_n_n432_ & new_n_n439_ & new_ni_4__;
  assign new_n_n108_ = new_n_n370_ & new_n_n110_ & new_n_n444_;
  assign new_n_n100_ = new_n_n212_ & new_n_n125_ & new_n_n277_;
  assign new_n_n92_ = new_n_n330_ & new_n_n96_ & new_n_n95_;
  assign new_n_n85_ = new_n_n319_ & new_n_n318_ & new_n_n371_;
  assign new_n_n457_ = ~new_ni_11__;
  assign new_n_n446_ = ~new_ni_50__;
  assign new_n_n430_ = ~new_ni_2__;
  assign new_n_n419_ = ~new_ni_34__;
  assign new_n_n408_ = ~new_ni_55__;
  assign new_n_n354_ = new_n_n439_ & new_n_n438_ & new_n_n437_;
  assign new_n_n339_ = new_n_n421_ & new_n_n420_ & new_n_n419_;
  assign new_n_n328_ = new_n_n340_ & new_n_n360_ & new_n_n387_;
  assign new_n_n318_ = new_n_n453_ & new_n_n436_ & new_n_n452_;
  assign new_n_n308_ = new_n_n434_ & new_n_n444_;
  assign new_n_n249_ = new_n_n252_ & new_n_n338_ & new_n_n266_;
  assign new_no_46__ = new_n_n240_ & new_n_n241_;
  assign new_n_n230_ = new_n_n429_ & new_n_n428_ & new_n_n438_;
  assign new_no_44__ = new_n_n220_ & new_n_n221_;
  assign new_n_n210_ = new_n_n271_ & new_n_n211_ & new_n_n286_;
  assign new_n_n162_ = new_n_n165_ & new_n_n194_ & new_n_n164_;
  assign new_n_n155_ = new_n_n419_ & new_n_n418_ & new_n_n417_;
  assign new_n_n145_ = new_n_n302_ & new_n_n301_ & new_n_n149_;
  assign new_n_n137_ = new_n_n426_ & new_ni_13__ & new_n_n456_;
  assign new_n_n127_ = new_n_n443_ & new_n_n421_ & new_ni_32__;
  assign new_no_26__ = new_n_n118_ & new_n_n117_ & new_n_n119_;
  assign new_n_n4_ = new_n_n387_ & new_n_n339_ & new_n_n293_;
  assign new_n_n456_ = ~new_ni_14__;
  assign new_n_n447_ = ~new_ni_46__;
  assign new_n_n429_ = ~new_ni_4__;
  assign new_n_n420_ = ~new_ni_33__;
  assign new_n_n398_ = ~new_ni_23__;
  assign new_no_59__ = new_n_n445_ & new_n_n363_;
  assign new_n_n338_ = new_n_n450_ & new_n_n449_ & new_n_n435_;
  assign new_n_n329_ = new_n_n343_ & new_n_n342_ & new_n_n341_;
  assign new_n_n317_ = new_ni_29__ & new_n_n443_ & new_ni_35__;
  assign new_n_n309_ = new_ni_55__ & new_n_n442_ & new_n_n445_;
  assign new_n_n248_ = new_n_n316_ & new_n_n278_ & new_n_n277_;
  assign new_n_n240_ = new_n_n273_ & new_n_n242_;
  assign new_n_n229_ = new_n_n437_ & new_n_n440_ & new_n_n427_;
  assign new_n_n220_ = new_n_n223_ & new_n_n222_ & new_n_n434_;
  assign new_n_n202_ = new_ni_54__ & new_n_n408_ & new_n_n442_;
  assign new_no_35__ = new_n_n163_ & new_n_n162_;
  assign new_n_n156_ = new_n_n424_ & new_n_n423_ & new_ni_21__;
  assign new_n_n144_ = new_n_n330_ & new_n_n148_ & new_n_n147_;
  assign new_no_28__ = new_n_n138_ & new_n_n139_;
  assign new_n_n126_ = new_n_n446_ & new_n_n412_ & new_n_n411_;
  assign new_n_n117_ = new_n_n122_ & new_n_n121_ & new_n_n120_;
  assign new_n_n5_ = new_n_n372_ & new_n_n294_ & new_n_n360_;
  assign new_n_n432_ = ~new_ni_0__;
  assign new_n_n421_ = ~new_ni_31__;
  assign new_n_n388_ = new_n_n392_ & new_n_n391_ & new_n_n390_;
  assign new_n_n371_ = new_ni_29__ & new_n_n443_ & new_n_n451_;
  assign new_n_n341_ = new_n_n425_ & new_n_n424_ & new_n_n423_;
  assign new_n_n330_ = new_n_n346_ & new_n_n345_ & new_n_n344_;
  assign new_n_n300_ = new_n_n412_ & new_n_n410_ & new_n_n409_;
  assign new_n_n290_ = new_n_n441_ & new_n_n414_ & new_n_n413_;
  assign new_n_n251_ = new_n_n268_ & new_n_n344_ & new_n_n395_;
  assign new_n_n241_ = new_n_n244_ & new_n_n236_ & new_n_n243_;
  assign new_n_n228_ = new_n_n455_ & new_n_n424_ & new_n_n423_;
  assign new_n_n212_ = new_n_n410_ & new_n_n409_ & new_n_n408_;
  assign new_n_n203_ = new_ni_29__ & new_n_n443_ & new_n_n420_;
  assign new_n_n164_ = new_n_n293_ & new_n_n168_ & new_n_n369_;
  assign new_no_32__ = new_n_n157_ & new_n_n142_;
  assign new_n_n143_ = new_n_n146_ & new_n_n145_ & new_n_n18_;
  assign new_n_n135_ = new_n_n343_ & new_n_n137_ & new_n_n185_;
  assign new_no_27__ = new_n_n130_ & new_n_n129_ & new_n_n131_;
  assign new_n_n118_ = new_n_n330_ & new_n_n181_ & new_n_n123_;
  assign new_n_n6_ = new_n_n268_ & new_n_n9_ & new_n_n8_;
  assign new_n_n431_ = ~new_ni_1__;
  assign new_n_n422_ = ~new_ni_21__;
  assign new_no_62__ = new_n_n382_ & new_n_n381_ & new_n_n444_;
  assign new_n_n380_ = new_ni_8__ & new_n_n458_ & new_n_n457_;
  assign new_n_n340_ = new_ni_20__ & new_n_n422_ & new_n_n433_;
  assign new_n_n331_ = new_n_n405_ & new_n_n434_ & new_n_n404_;
  assign new_n_n299_ = new_n_n405_ & new_n_n434_ & new_ni_63__;
  assign new_n_n291_ = new_n_n448_ & new_n_n415_ & new_n_n447_;
  assign new_n_n250_ = new_n_n253_ & new_n_n352_ & new_n_n351_;
  assign new_n_n242_ = new_n_n369_ & new_n_n167_ & new_n_n332_;
  assign new_n_n219_ = new_n_n432_ & new_ni_1__ & new_n_n430_;
  assign new_n_n211_ = new_n_n213_ & new_n_n212_ & new_n_n264_;
  assign new_no_41__ = new_n_n204_ & new_n_n205_;
  assign new_n_n163_ = new_n_n167_ & new_n_n166_ & new_n_n434_;
  assign new_n_n157_ = new_ni_46__ & new_n_n446_ & new_n_n445_;
  assign new_no_30__ = new_n_n144_ & new_n_n143_ & new_n_n285_;
  assign new_n_n136_ = new_n_n412_ & new_n_n411_ & new_n_n410_;
  assign new_n_n128_ = new_n_n423_ & new_n_n401_ & new_n_n422_;
  assign new_n_n119_ = new_n_n124_ & new_n_n277_;
  assign new_n_n7_ = new_n_n448_ & new_ni_45__ & new_n_n447_;
  assign new_n_n453_ = ~new_ni_25__;
  assign new_n_n442_ = ~new_ni_56__;
  assign new_n_n412_ = ~new_ni_51__;
  assign new_n_n401_ = ~new_ni_20__;
  assign new_n_n390_ = new_n_n444_ & new_n_n445_;
  assign new_n_n381_ = new_n_n392_ & new_n_n384_ & new_n_n383_;
  assign new_n_n379_ = new_n_n453_ & new_n_n452_ & new_ni_29__;
  assign new_n_n369_ = new_n_n447_ & new_n_n441_ & new_n_n446_;
  assign new_n_n360_ = new_n_n454_ & new_n_n453_ & new_n_n436_;
  assign new_n_n350_ = new_n_n354_ & new_n_n362_ & new_n_n353_;
  assign new_no_56__ = new_n_n323_ & new_n_n322_ & new_n_n324_;
  assign new_n_n311_ = new_n_n315_ & new_n_n314_ & new_n_n313_;
  assign new_n_n302_ = new_n_n415_ & new_n_n447_ & new_n_n441_;
  assign new_n_n292_ = new_n_n449_ & new_n_n435_ & new_n_n416_;
  assign new_n_n289_ = new_n_n446_ & new_n_n412_ & new_n_n410_;
  assign new_n_n279_ = new_ni_48__ & new_n_n413_ & new_n_n446_;
  assign new_n_n269_ = new_n_n271_ & new_n_n270_ & new_n_n199_;
  assign new_no_49__ = new_n_n260_ & new_n_n198_;
  assign new_no_47__ = new_n_n246_ & new_n_n247_;
  assign new_n_n233_ = new_n_n263_ & new_n_n236_ & new_n_n235_;
  assign new_n_n223_ = new_n_n338_ & new_n_n337_ & new_n_n369_;
  assign new_no_43__ = new_n_n214_ & new_n_n215_;
  assign new_n_n204_ = new_n_n206_ & new_n_n207_;
  assign new_n_n192_ = new_n_n237_ & new_n_n368_ & new_n_n273_;
  assign new_n_n183_ = new_n_n400_ & new_n_n420_ & new_n_n419_;
  assign new_n_n173_ = new_n_n444_ & new_ni_61__ & new_n_n434_;
  assign new_n_n160_ = new_ni_39__ & new_n_n449_ & new_n_n448_;
  assign new_n_n151_ = new_n_n146_ & new_n_n153_ & new_n_n28_;
  assign new_n_n149_ = new_n_n412_ & new_ni_52__ & new_n_n410_;
  assign new_n_n140_ = new_ni_25__ & new_n_n452_ & new_ni_29__;
  assign new_n_n130_ = new_n_n330_ & new_n_n135_ & new_n_n123_;
  assign new_n_n120_ = new_n_n126_ & new_n_n212_ & new_n_n125_;
  assign new_n_n98_ = new_n_n102_ & new_n_n101_ & new_n_n100_;
  assign new_n_n89_ = new_n_n90_ & new_n_n320_ & new_n_n372_;
  assign new_n_n0_ = new_n_n2_ & new_n_n3_;
  assign new_n_n452_ = ~new_ni_28__;
  assign new_n_n443_ = ~new_ni_30__;
  assign new_n_n411_ = ~new_ni_52__;
  assign new_n_n402_ = ~new_ni_13__;
  assign new_n_n389_ = new_n_n395_ & new_n_n394_ & new_n_n393_;
  assign new_n_n382_ = new_n_n395_ & new_n_n394_ & new_n_n387_;
  assign new_n_n378_ = new_n_n443_ & new_n_n451_ & new_n_n450_;
  assign new_n_n370_ = new_n_n450_ & new_n_n449_ & new_n_n448_;
  assign new_n_n359_ = new_n_n435_ & new_n_n448_ & new_n_n447_;
  assign new_n_n351_ = new_n_n436_ & new_n_n452_ & new_ni_29__;
  assign new_n_n321_ = new_n_n432_ & new_n_n439_ & new_n_n438_;
  assign new_n_n312_ = new_n_n434_ & new_n_n368_;
  assign new_n_n301_ = new_n_n414_ & new_n_n413_ & new_n_n446_;
  assign new_n_n293_ = new_n_n418_ & new_n_n451_ & new_n_n450_;
  assign new_n_n288_ = new_n_n409_ & new_n_n408_ & new_n_n442_;
  assign new_no_52__ = new_n_n280_ & new_n_n281_;
  assign new_no_50__ = new_n_n269_ & new_n_n297_;
  assign new_n_n260_ = new_n_n261_ & new_n_n262_;
  assign new_n_n237_ = new_n_n446_ & new_n_n412_ & new_n_n408_;
  assign new_n_n232_ = new_n_n286_ & new_n_n234_;
  assign new_n_n224_ = new_n_n351_ & new_n_n227_ & new_n_n267_;
  assign new_n_n213_ = new_ni_49__ & new_n_n446_ & new_n_n412_;
  assign new_n_n205_ = new_n_n263_ & new_n_n236_ & new_n_n208_;
  assign new_n_n201_ = new_n_n203_ & new_n_n267_ & new_n_n338_;
  assign new_n_n182_ = new_n_n418_ & new_n_n417_ & new_n_n451_;
  assign new_no_37__ = new_n_n175_ & new_n_n174_ & new_n_n176_;
  assign new_n_n159_ = new_n_n445_ & new_n_n446_;
  assign new_n_n152_ = new_n_n330_ & new_n_n154_ & new_n_n147_;
  assign new_n_n148_ = new_n_n343_ & new_n_n342_ & new_n_n150_;
  assign new_no_29__ = new_n_n141_ & new_n_n142_;
  assign new_n_n129_ = new_n_n134_ & new_n_n133_ & new_n_n132_;
  assign new_n_n121_ = new_n_n292_ & new_n_n291_ & new_n_n290_;
  assign new_no_23__ = new_n_n99_ & new_n_n98_ & new_n_n124_;
  assign new_n_n90_ = new_ni_0__ & new_n_n439_ & new_n_n438_;
  assign new_n_n1_ = new_n_n6_ & new_n_n5_ & new_n_n4_;
  assign new_n_n455_ = ~new_ni_15__;
  assign new_n_n444_ = ~new_ni_60__;
  assign new_n_n428_ = ~new_ni_5__;
  assign new_n_n410_ = ~new_ni_53__;
  assign new_n_n399_ = ~new_ni_19__;
  assign new_n_n392_ = new_n_n451_ & new_n_n450_ & new_n_n449_;
  assign new_n_n383_ = new_n_n446_ & new_n_n442_ & new_n_n445_;
  assign new_n_n377_ = new_n_n449_ & new_n_n448_ & new_n_n447_;
  assign new_n_n367_ = new_n_n373_ & new_n_n372_ & new_n_n78_;
  assign new_n_n362_ = new_n_n440_ & new_n_n458_ & new_n_n457_;
  assign new_n_n352_ = new_n_n433_ & new_n_n454_ & new_n_n453_;
  assign new_n_n337_ = new_n_n416_ & new_n_n448_ & new_n_n415_;
  assign new_n_n326_ = new_n_n337_ & new_n_n336_ & new_n_n335_;
  assign new_n_n320_ = new_n_n437_ & new_n_n440_ & new_n_n458_;
  assign new_n_n310_ = new_ni_29__ & new_n_n443_ & new_n_n418_;
  assign new_n_n304_ = new_n_n420_ & new_n_n419_ & new_n_n418_;
  assign new_n_n294_ = new_n_n424_ & new_n_n423_ & new_n_n433_;
  assign new_n_n287_ = new_n_n407_ & new_n_n445_ & new_n_n406_;
  assign new_n_n277_ = new_n_n406_ & new_n_n444_ & new_n_n405_;
  assign new_n_n271_ = new_n_n392_ & new_n_n303_ & new_n_n302_;
  assign new_n_n261_ = new_n_n286_ & new_n_n264_;
  assign new_n_n247_ = new_n_n251_ & new_n_n250_ & new_n_n249_;
  assign new_n_n238_ = new_n_n448_ & new_n_n447_ & new_n_n441_;
  assign new_no_45__ = new_n_n232_ & new_n_n233_;
  assign new_n_n221_ = new_n_n226_ & new_n_n225_ & new_n_n224_;
  assign new_n_n215_ = new_n_n218_ & new_n_n217_ & new_n_n272_;
  assign new_n_n206_ = new_n_n434_ & new_n_n277_;
  assign new_n_n200_ = new_n_n266_ & new_n_n316_ & new_n_n202_;
  assign new_no_39__ = new_n_n192_ & new_n_n191_;
  assign new_n_n174_ = new_n_n179_ & new_n_n178_ & new_n_n177_;
  assign new_n_n161_ = new_n_n456_ & new_n_n455_ & new_n_n452_;
  assign new_n_n153_ = new_n_n302_ & new_n_n301_ & new_n_n300_;
  assign new_n_n147_ = new_n_n352_ & new_n_n351_ & new_n_n227_;
  assign new_n_n138_ = new_n_n390_ & new_n_n391_;
  assign new_n_n132_ = new_n_n136_ & new_n_n288_ & new_n_n287_;
  assign new_n_n122_ = new_n_n127_ & new_n_n304_ & new_n_n105_;
  assign new_n_n116_ = new_ni_24__ & new_n_n453_ & new_n_n452_;
  assign new_n_n107_ = new_ni_16__ & new_n_n424_ & new_n_n423_;
  assign new_n_n2_ = new_n_n212_ & new_n_n264_ & new_n_n286_;
  assign new_n_n454_ = ~new_ni_24__;
  assign new_n_n445_ = ~new_ni_58__;
  assign new_n_n418_ = ~new_ni_35__;
  assign new_n_n409_ = ~new_ni_54__;
  assign new_n_n400_ = ~new_ni_32__;
  assign new_n_n391_ = new_n_n448_ & new_n_n447_ & new_n_n446_;
  assign new_n_n384_ = new_n_n448_ & new_n_n447_ & new_ni_47__;
  assign new_n_n376_ = new_n_n441_ & new_n_n446_ & new_n_n442_;
  assign new_n_n368_ = new_n_n442_ & new_n_n445_ & new_n_n444_;
  assign new_n_n361_ = new_n_n456_ & new_n_n455_ & new_ni_22__;
  assign new_n_n353_ = new_n_n456_ & new_n_n455_ & new_ni_18__;
  assign new_n_n336_ = new_n_n447_ & new_n_n441_ & new_n_n414_;
  assign new_n_n327_ = new_n_n339_ & new_n_n182_ & new_n_n338_;
  assign new_n_n319_ = new_n_n423_ & new_n_n433_ & new_n_n454_;
  assign new_no_55__ = new_n_n312_ & new_n_n311_;
  assign new_n_n303_ = new_n_n435_ & new_n_n416_ & new_n_n448_;
  assign new_n_n295_ = new_ni_12__ & new_n_n456_ & new_n_n455_;
  assign new_n_n286_ = new_n_n444_ & new_n_n405_ & new_n_n434_;
  assign new_n_n278_ = new_n_n408_ & new_n_n442_ & new_n_n445_;
  assign new_n_n270_ = new_n_n301_ & new_n_n300_ & new_n_n274_;
  assign new_n_n262_ = new_n_n266_ & new_n_n316_ & new_n_n265_;
  assign new_n_n246_ = new_n_n434_ & new_n_n248_;
  assign new_n_n239_ = new_ni_29__ & new_n_n443_ & new_ni_34__;
  assign new_n_n231_ = new_n_n432_ & new_ni_2__ & new_n_n439_;
  assign new_n_n222_ = new_n_n300_ & new_n_n278_ & new_n_n277_;
  assign new_n_n214_ = new_n_n271_ & new_n_n216_ & new_n_n273_;
  assign new_n_n207_ = new_n_n266_ & new_n_n316_ & new_n_n278_;
  assign new_n_n199_ = new_n_n273_ & new_n_n332_;
  assign new_n_n191_ = new_n_n251_ & new_n_n194_ & new_n_n193_;
  assign new_n_n184_ = new_n_n423_ & new_ni_19__ & new_n_n401_;
  assign new_no_34__ = new_n_n161_ & new_n_n34_ & new_ni_58__;
  assign new_n_n154_ = new_n_n343_ & new_n_n342_ & new_n_n156_;
  assign new_n_n146_ = new_n_n155_ & new_n_n392_ & new_n_n303_;
  assign new_n_n139_ = new_n_n366_ & new_n_n140_ & new_n_n392_;
  assign new_n_n131_ = new_n_n285_ & new_n_n286_;
  assign new_n_n123_ = new_n_n128_ & new_n_n352_ & new_n_n351_;
  assign new_n_n115_ = new_ni_29__ & new_n_n451_ & new_n_n450_;
  assign new_no_24__ = new_n_n108_ & new_n_n109_;
  assign new_n_n3_ = new_n_n292_ & new_n_n7_ & new_n_n316_;
  assign new_n_n78_ = new_n_n454_ & new_n_n453_ & new_n_n452_;
  assign new_n_n69_ = new_n_n70_ & new_n_n378_ & new_n_n377_;
  assign new_n_n61_ = new_n_n351_ & new_n_n378_ & new_n_n63_;
  assign new_n_n53_ = new_n_n423_ & new_n_n399_ & new_n_n401_;
  assign new_n_n43_ = new_n_n451_ & new_ni_38__ & new_n_n450_;
  assign new_no_19__ = new_n_n79_ & new_n_n297_;
  assign new_n_n68_ = new_n_n358_ & new_n_n376_;
  assign new_n_n62_ = new_n_n64_ & new_n_n395_ & new_n_n394_;
  assign new_n_n52_ = new_n_n422_ & new_n_n433_ & new_ni_23__;
  assign new_n_n44_ = new_n_n422_ & new_n_n433_ & new_n_n398_;
  assign new_n_n79_ = new_n_n271_ & new_n_n81_ & new_n_n80_;
  assign new_no_16__ = new_n_n62_ & new_n_n69_ & new_n_n68_;
  assign new_no_13__ = new_n_n62_ & new_n_n61_ & new_n_n60_;
  assign new_n_n54_ = new_n_n455_ & new_ni_28__ & new_ni_29__;
  assign new_no_9__ = new_n_n46_ & new_n_n45_ & new_n_n47_;
  assign new_n_n80_ = new_n_n82_ & new_n_n332_;
  assign new_n_n67_ = new_ni_10__ & new_n_n456_ & new_n_n455_;
  assign new_n_n60_ = new_n_n369_ & new_n_n368_ & new_n_n434_;
  assign new_no_10__ = new_n_n451_ & new_n_n54_;
  assign new_n_n45_ = new_n_n49_ & new_n_n271_ & new_n_n48_;
  assign new_no_0__ = new_n_n0_ & new_n_n1_;
  assign new_n_n81_ = new_n_n301_ & new_n_n300_ & new_n_n333_;
  assign new_n_n37_ = new_n_n455_ & new_n_n452_ & new_ni_29__;
  assign new_n_n28_ = new_n_n333_ & new_n_n332_ & new_n_n331_;
  assign new_n_n18_ = new_n_n288_ & new_n_n287_ & new_n_n286_;
  assign new_n_n9_ = new_n_n428_ & new_n_n438_ & new_n_n437_;
  assign new_n_n82_ = new_n_n405_ & new_n_n434_ & new_ni_64__;
  assign new_n_n36_ = new_ni_43__ & new_n_n451_;
  assign new_n_n29_ = new_n_n336_ & new_n_n335_ & new_n_n334_;
  assign new_n_n17_ = new_n_n21_ & new_n_n20_ & new_n_n19_;
  assign new_no_1__ = new_n_n10_ & new_n_n11_;
  assign new_no_7__ = new_n_n36_ & new_n_n37_;
  assign new_n_n26_ = new_n_n403_ & new_n_n28_;
  assign new_n_n20_ = new_n_n23_ & new_n_n338_ & new_n_n22_;
  assign new_n_n10_ = new_n_n12_ & new_n_n13_;
  assign new_n_n35_ = new_ni_14__ & new_n_n455_ & new_n_n452_;
  assign new_n_n27_ = new_n_n49_ & new_n_n30_ & new_n_n29_;
  assign new_n_n19_ = new_n_n302_ & new_n_n301_ & new_n_n136_;
  assign new_n_n11_ = new_n_n14_ & new_n_n5_ & new_n_n4_;
  assign new_n_n59_ = new_n_n439_ & new_ni_6__ & new_n_n437_;
  assign new_n_n50_ = new_n_n53_ & new_n_n52_ & new_n_n360_;
  assign new_n_n40_ = new_n_n125_ & new_n_n277_ & new_n_n124_;
  assign new_n_n32_ = new_n_n448_ & new_ni_44__ & new_n_n415_;
  assign new_n_n22_ = new_n_n416_ & new_n_n448_ & new_n_n396_;
  assign new_n_n12_ = new_n_n288_ & new_n_n332_ & new_n_n273_;
  assign new_n_n58_ = new_n_n456_ & new_n_n455_ & new_n_n454_;
  assign new_n_n51_ = new_n_n421_ & new_n_n400_ & new_n_n420_;
  assign new_n_n39_ = new_n_n330_ & new_n_n181_ & new_n_n31_;
  assign new_n_n33_ = new_n_n451_ & new_n_n397_ & new_n_n450_;
  assign new_n_n21_ = new_n_n25_ & new_n_n24_ & new_n_n304_;
  assign new_n_n13_ = new_n_n292_ & new_n_n238_ & new_n_n289_;
  assign new_n_n74_ = new_ni_3__ & new_n_n437_ & new_n_n440_;
  assign new_no_15__ = new_n_n67_ & new_n_n365_ & new_n_n66_;
  assign new_n_n38_ = new_n_n49_ & new_n_n42_ & new_n_n41_;
  assign new_n_n30_ = new_n_n33_ & new_n_n292_ & new_n_n32_;
  assign new_n_n24_ = new_n_n443_ & new_n_n421_ & new_n_n400_;
  assign new_n_n14_ = new_n_n268_ & new_n_n15_ & new_n_n8_;
  assign new_n_n73_ = new_n_n74_ & new_n_n395_ & new_n_n394_;
  assign new_n_n66_ = new_n_n445_ & new_n_n448_;
  assign new_no_8__ = new_n_n39_ & new_n_n38_ & new_n_n40_;
  assign new_n_n31_ = new_n_n53_ & new_n_n44_ & new_n_n360_;
  assign new_n_n23_ = new_n_n417_ & new_n_n451_ & new_n_n397_;
  assign new_n_n15_ = new_ni_5__ & new_n_n438_ & new_n_n437_;
  assign new_no_18__ = new_n_n77_ & new_n_n76_ & new_n_n75_;
  assign new_n_n72_ = new_n_n387_ & new_n_n392_ & new_n_n238_;
  assign new_no_14__ = new_n_n366_ & new_n_n365_ & new_n_n65_;
  assign new_n_n55_ = new_n_n238_ & new_n_n383_ & new_n_n308_;
  assign new_n_n46_ = new_n_n330_ & new_n_n181_ & new_n_n50_;
  assign new_no_3__ = new_n_n39_ & new_n_n27_ & new_n_n26_;
  assign new_no_2__ = new_n_n39_ & new_n_n17_ & new_n_n16_;
  assign new_n_n75_ = new_ni_62__ & new_n_n368_;
  assign new_n_n71_ = new_n_n308_ & new_n_n383_;
  assign new_n_n65_ = new_n_n448_ & new_ni_50__ & new_n_n445_;
  assign new_no_12__ = new_n_n57_ & new_n_n56_ & new_n_n55_;
  assign new_n_n47_ = new_n_n287_ & new_n_n286_ & new_n_n285_;
  assign new_n_n25_ = new_ni_27__ & new_n_n452_ & new_ni_29__;
  assign new_n_n16_ = new_n_n285_ & new_n_n18_;
  assign new_n_n76_ = new_n_n371_ & new_n_n370_ & new_n_n369_;
  assign new_no_17__ = new_n_n73_ & new_n_n72_ & new_n_n71_;
  assign new_n_n63_ = new_n_n449_ & new_ni_41__ & new_n_n448_;
  assign new_n_n57_ = new_n_n59_ & new_n_n362_ & new_n_n58_;
  assign new_n_n48_ = new_n_n301_ & new_n_n136_ & new_n_n288_;
  assign new_n_n42_ = new_n_n43_ & new_n_n292_ & new_n_n291_;
  assign new_no_6__ = new_n_n34_ & new_n_n35_;
  assign new_n_n77_ = new_n_n320_ & new_n_n372_ & new_n_n78_;
  assign new_n_n70_ = new_ni_26__ & new_n_n452_ & new_ni_29__;
  assign new_n_n64_ = new_n_n439_ & new_n_n437_ & new_n_n440_;
  assign new_n_n56_ = new_n_n318_ & new_n_n371_ & new_n_n338_;
  assign new_n_n49_ = new_n_n387_ & new_n_n51_ & new_n_n155_;
  assign new_n_n41_ = new_n_n290_ & new_n_n126_ & new_n_n212_;
  assign new_n_n34_ = new_ni_29__ & new_n_n451_ & new_n_n448_;
endmodule


