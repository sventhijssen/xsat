// Benchmark "top" written by ABC on Fri Mar 31 12:08:35 2023

module top ( 
    pv16_9_, pv40_15_, pv88_6_, pv28_10_, pv88_7_, pv109_1_, pv118_3_,
    pv2_0_, pv40_13_, pv52_10_, pv109_2_, pv128_3_, pv2_1_, pv40_14_,
    pv52_11_, pv88_9_, pv109_3_, pv16_5_, pv40_11_, pv76_3_, pv88_2_,
    pv88_15_, pv100_14_, pv128_1_, pv16_13_, pv52_13_, pv76_2_, pv88_3_,
    pv100_13_, pv128_2_, pv16_7_, pv16_14_, pv52_14_, pv76_1_, pv88_13_,
    pv118_2_, pv16_6_, pv16_15_, pv40_10_, pv52_15_, pv88_5_, pv88_14_,
    pv100_15_, pv118_1_, pv128_0_, pv4_0_, pv52_9_, pv88_11_, pv100_3_,
    pv100_10_, pv121_2_, pv132_0_, pv4_1_, pv28_9_, pv64_1_, pv121_3_,
    pv16_10_, pv28_6_, pv100_5_, pv16_11_, pv28_7_, pv88_10_, pv100_6_,
    pv100_11_, pv121_1_, pv76_14_, pv28_5_, pv64_5_, pv76_15_, pv28_2_,
    pv64_2_, pv100_1_, pv28_3_, pv64_3_, pv100_2_, pv52_1_, pv76_10_,
    pv103_2_, pv124_1_, pv28_1_, pv64_9_, pv76_11_, pv103_3_, pv124_2_,
    pv52_3_, pv64_6_, pv64_15_, pv52_2_, pv64_7_, pv76_13_, pv52_5_,
    pv100_7_, pv112_2_, pv112_1_, pv132_3_, pv133_0_, pv52_7_, pv100_9_,
    pv132_2_, pv40_1_, pv52_6_, pv103_1_, pv112_3_, pv132_1_, pv16_1_,
    pv40_2_, pv76_7_, pv106_1_, pv40_3_, pv64_10_, pv76_6_, pv106_2_,
    pv16_3_, pv28_15_, pv76_5_, pv106_3_, pv16_2_, pv40_5_, pv88_1_,
    pv28_13_, pv40_6_, pv64_13_, pv115_1_, pv28_14_, pv40_7_, pv64_14_,
    pv28_11_, pv64_11_, pv76_9_, pv115_3_, pv124_3_, pv40_9_, pv115_2_,
    pv167_11_, pv199_9_, pv167_12_, pv199_8_, pv167_13_, pv167_14_,
    pv151_1_, pv199_5_, pv151_0_, pv183_10_, pv199_4_, pv151_3_, pv183_11_,
    pv199_7_, pv151_2_, pv167_10_, pv183_12_, pv199_6_, pv167_4_, pv199_1_,
    pv167_5_, pv199_0_, pv167_2_, pv199_3_, pv167_3_, pv199_2_, pv167_8_,
    pv199_14_, pv167_9_, pv199_15_, pv167_6_, pv199_12_, pv167_7_,
    pv199_13_, pv199_10_, pv199_11_, pv167_0_, pv183_6_, pv167_1_,
    pv183_7_, pv183_8_, pv183_9_, pv151_5_, pv151_14_, pv183_2_, pv183_13_,
    pv151_4_, pv151_15_, pv183_3_, pv183_14_, pv151_7_, pv151_12_,
    pv183_4_, pv183_15_, pv151_6_, pv151_13_, pv183_5_, pv151_9_,
    pv151_10_, pv167_15_, pv151_8_, pv151_11_, pv135_1_, pv183_0_,
    pv135_0_, pv183_1_  );
  input  pv16_9_, pv40_15_, pv88_6_, pv28_10_, pv88_7_, pv109_1_,
    pv118_3_, pv2_0_, pv40_13_, pv52_10_, pv109_2_, pv128_3_, pv2_1_,
    pv40_14_, pv52_11_, pv88_9_, pv109_3_, pv16_5_, pv40_11_, pv76_3_,
    pv88_2_, pv88_15_, pv100_14_, pv128_1_, pv16_13_, pv52_13_, pv76_2_,
    pv88_3_, pv100_13_, pv128_2_, pv16_7_, pv16_14_, pv52_14_, pv76_1_,
    pv88_13_, pv118_2_, pv16_6_, pv16_15_, pv40_10_, pv52_15_, pv88_5_,
    pv88_14_, pv100_15_, pv118_1_, pv128_0_, pv4_0_, pv52_9_, pv88_11_,
    pv100_3_, pv100_10_, pv121_2_, pv132_0_, pv4_1_, pv28_9_, pv64_1_,
    pv121_3_, pv16_10_, pv28_6_, pv100_5_, pv16_11_, pv28_7_, pv88_10_,
    pv100_6_, pv100_11_, pv121_1_, pv76_14_, pv28_5_, pv64_5_, pv76_15_,
    pv28_2_, pv64_2_, pv100_1_, pv28_3_, pv64_3_, pv100_2_, pv52_1_,
    pv76_10_, pv103_2_, pv124_1_, pv28_1_, pv64_9_, pv76_11_, pv103_3_,
    pv124_2_, pv52_3_, pv64_6_, pv64_15_, pv52_2_, pv64_7_, pv76_13_,
    pv52_5_, pv100_7_, pv112_2_, pv112_1_, pv132_3_, pv133_0_, pv52_7_,
    pv100_9_, pv132_2_, pv40_1_, pv52_6_, pv103_1_, pv112_3_, pv132_1_,
    pv16_1_, pv40_2_, pv76_7_, pv106_1_, pv40_3_, pv64_10_, pv76_6_,
    pv106_2_, pv16_3_, pv28_15_, pv76_5_, pv106_3_, pv16_2_, pv40_5_,
    pv88_1_, pv28_13_, pv40_6_, pv64_13_, pv115_1_, pv28_14_, pv40_7_,
    pv64_14_, pv28_11_, pv64_11_, pv76_9_, pv115_3_, pv124_3_, pv40_9_,
    pv115_2_;
  output pv167_11_, pv199_9_, pv167_12_, pv199_8_, pv167_13_, pv167_14_,
    pv151_1_, pv199_5_, pv151_0_, pv183_10_, pv199_4_, pv151_3_, pv183_11_,
    pv199_7_, pv151_2_, pv167_10_, pv183_12_, pv199_6_, pv167_4_, pv199_1_,
    pv167_5_, pv199_0_, pv167_2_, pv199_3_, pv167_3_, pv199_2_, pv167_8_,
    pv199_14_, pv167_9_, pv199_15_, pv167_6_, pv199_12_, pv167_7_,
    pv199_13_, pv199_10_, pv199_11_, pv167_0_, pv183_6_, pv167_1_,
    pv183_7_, pv183_8_, pv183_9_, pv151_5_, pv151_14_, pv183_2_, pv183_13_,
    pv151_4_, pv151_15_, pv183_3_, pv183_14_, pv151_7_, pv151_12_,
    pv183_4_, pv183_15_, pv151_6_, pv151_13_, pv183_5_, pv151_9_,
    pv151_10_, pv167_15_, pv151_8_, pv151_11_, pv135_1_, pv183_0_,
    pv135_0_, pv183_1_;
  wire new_n_n174_, new_n_n154_, new_n_n118_, new_n_n184_, new_n_n116_,
    new_n_n78_, new_n_n85_, new_n_n197_, new_n_n149_, new_n_n160_,
    new_n_n93_, new_n_n70_, new_n_n199_, new_n_n156_, new_n_n158_,
    new_n_n101_, new_n_n91_, new_n_n175_, new_n_n159_, new_n_n144_,
    new_n_n123_, new_n_n106_, new_n_n107_, new_n_n74_, new_n_n173_,
    new_n_n157_, new_n_n146_, new_n_n121_, new_n_n109_, new_n_n72_,
    new_n_n188_, new_n_n180_, new_n_n155_, new_n_n148_, new_n_n100_,
    new_n_n87_, new_n_n190_, new_n_n178_, new_n_n161_, new_n_n153_,
    new_n_n102_, new_n_n108_, new_n_n104_, new_n_n89_, new_n_n68_,
    new_n_n200_, new_n_n162_, new_n_n111_, new_n_n120_, new_n_n112_,
    new_n_n83_, new_n_n75_, new_n_n198_, new_n_n186_, new_n_n128_,
    new_n_n81_, new_n_n185_, new_n_n189_, new_n_n119_, new_n_n183_,
    new_n_n187_, new_n_n113_, new_n_n117_, new_n_n110_, new_n_n76_,
    new_n_n131_, new_n_n191_, new_n_n127_, new_n_n129_, new_n_n194_,
    new_n_n147_, new_n_n124_, new_n_n192_, new_n_n145_, new_n_n122_,
    new_n_n172_, new_n_n136_, new_n_n98_, new_n_n84_, new_n_n196_,
    new_n_n126_, new_n_n134_, new_n_n96_, new_n_n82_, new_n_n168_,
    new_n_n142_, new_n_n130_, new_n_n170_, new_n_n140_, new_n_n133_,
    new_n_n167_, new_n_n115_, new_n_n92_, new_n_n94_, new_n_n69_,
    new_n_n105_, new_n_n163_, new_n_n114_, new_n_n71_, new_n_n152_,
    new_n_n165_, new_n_n79_, new_n_n90_, new_n_n73_, new_n_n176_,
    new_n_n171_, new_n_n139_, new_n_n99_, new_n_n169_, new_n_n137_,
    new_n_n141_, new_n_n97_, new_n_n193_, new_n_n177_, new_n_n143_,
    new_n_n95_, new_n_n195_, new_n_n151_, new_n_n103_, new_n_n181_,
    new_n_n166_, new_n_n125_, new_n_n77_, new_n_n179_, new_n_n164_,
    new_n_n132_, new_n_n182_, new_n_n135_, new_n_n138_, new_n_n86_,
    new_n_n80_, new_n_n150_, new_n_n88_, new_n_n55_, new_nv236_,
    new_nv247_, new_n_n46_, new_nv257_, new_nv268_, new_n_n54_, new_nv235_,
    new_nv248_, new_n_n47_, new_nv258_, new_nv267_, new_nv217_, new_n_n64_,
    new_nv249_, new_n_n44_, new_nv255_, new_nv266_, new_nv218_, new_n_n65_,
    new_nv250_, new_n_n45_, new_nv256_, new_nv265_, new_nv208_, new_n_n53_,
    new_n_n42_, new_nv261_, new_nv272_, new_nv327_, new_nv200_, new_nv207_,
    new_n_n52_, new_n_n43_, new_nv262_, new_nv271_, new_n_n51_, new_nv252_,
    new_nv259_, new_nv270_, new_n_n50_, new_nv251_, new_nv260_, new_nv269_,
    new_n_n67_, new_nv212_, new_nv223_, new_n_n58_, new_nv233_, new_nv244_,
    new_nv331_, new_n_n66_, new_nv211_, new_nv224_, new_n_n59_, new_nv234_,
    new_nv243_, new_nv330_, new_nv201_, new_nv210_, new_nv225_, new_n_n56_,
    new_nv231_, new_nv242_, new_nv329_, new_nv202_, new_nv209_, new_nv226_,
    new_n_n57_, new_nv232_, new_nv241_, new_nv328_, new_nv205_, new_nv216_,
    new_nv219_, new_n_n62_, new_nv229_, new_nv240_, new_nv253_, new_nv264_,
    new_n_n3_, new_nv206_, new_nv215_, new_nv220_, new_n_n63_, new_nv230_,
    new_nv239_, new_nv254_, new_nv263_, new_n_n4_, new_nv203_, new_nv214_,
    new_nv221_, new_n_n60_, new_nv227_, new_nv238_, new_nv245_, new_n_n48_,
    new_n_n5_, new_nv204_, new_nv213_, new_nv222_, new_n_n61_, new_nv228_,
    new_nv237_, new_nv246_, new_n_n49_, new_nv332_, new_n_n38_, new_nv277_,
    new_nv288_, new_n_n29_, new_n_n18_, new_n_n39_, new_nv278_, new_nv287_,
    new_n_n28_, new_n_n19_, new_n_n40_, new_nv279_, new_nv290_, new_nv297_,
    new_n_n20_, new_n_n41_, new_nv280_, new_nv289_, new_nv298_, new_n_n21_,
    new_n_n2_, new_nv274_, new_nv305_, new_nv316_, new_n_n13_, new_nv326_,
    new_nv273_, new_nv306_, new_nv315_, new_n_n12_, new_nv325_, new_nv307_,
    new_nv318_, new_n_n15_, new_nv324_, new_nv308_, new_nv317_, new_n_n14_,
    new_nv323_, new_nv291_, new_n_n26_, new_nv301_, new_nv312_, new_n_n17_,
    new_n_n6_, new_nv292_, new_n_n27_, new_nv302_, new_nv311_, new_n_n16_,
    new_n_n7_, new_n_n33_, new_nv282_, new_nv303_, new_nv314_, new_nv321_,
    new_n_n8_, new_n_n32_, new_nv281_, new_nv304_, new_nv313_, new_nv322_,
    new_n_n9_, new_n_n34_, new_n_n31_, new_nv284_, new_nv295_, new_n_n22_,
    new_nv319_, new_n_n10_, new_n_n35_, new_n_n30_, new_nv283_, new_nv296_,
    new_n_n23_, new_nv320_, new_n_n11_, new_n_n36_, new_nv275_, new_nv286_,
    new_nv293_, new_n_n24_, new_nv299_, new_nv310_, new_n_n37_, new_nv276_,
    new_nv285_, new_nv294_, new_n_n25_, new_nv300_, new_nv309_;
  assign new_n_n174_ = pv16_9_;
  assign new_n_n154_ = pv40_15_;
  assign new_n_n118_ = pv88_6_;
  assign pv167_11_ = new_n_n45_;
  assign pv199_9_ = new_n_n23_;
  assign new_n_n184_ = pv28_10_;
  assign new_n_n116_ = pv88_7_;
  assign new_n_n78_ = pv109_1_;
  assign new_n_n85_ = pv118_3_;
  assign pv167_12_ = new_n_n12_;
  assign pv199_8_ = new_n_n7_;
  assign new_n_n197_ = pv2_0_;
  assign new_n_n149_ = pv40_13_;
  assign new_n_n160_ = pv52_10_;
  assign new_n_n93_ = pv109_2_;
  assign new_n_n70_ = pv128_3_;
  assign pv167_13_ = new_n_n44_;
  assign new_n_n199_ = pv2_1_;
  assign new_n_n156_ = pv40_14_;
  assign new_n_n158_ = pv52_11_;
  assign new_n_n101_ = pv88_9_;
  assign new_n_n91_ = pv109_3_;
  assign pv167_14_ = new_n_n43_;
  assign new_n_n175_ = pv16_5_;
  assign new_n_n159_ = pv40_11_;
  assign new_n_n144_ = pv76_3_;
  assign new_n_n123_ = pv88_2_;
  assign new_n_n106_ = pv88_15_;
  assign new_n_n107_ = pv100_14_;
  assign new_n_n74_ = pv128_1_;
  assign pv151_1_ = new_n_n65_;
  assign pv199_5_ = new_n_n26_;
  assign new_n_n173_ = pv16_13_;
  assign new_n_n157_ = pv52_13_;
  assign new_n_n146_ = pv76_2_;
  assign new_n_n121_ = pv88_3_;
  assign new_n_n109_ = pv100_13_;
  assign new_n_n72_ = pv128_2_;
  assign pv151_0_ = new_n_n5_;
  assign pv183_10_ = new_n_n34_;
  assign pv199_4_ = new_n_n8_;
  assign new_n_n188_ = pv16_7_;
  assign new_n_n180_ = pv16_14_;
  assign new_n_n155_ = pv52_14_;
  assign new_n_n148_ = pv76_1_;
  assign new_n_n100_ = pv88_13_;
  assign new_n_n87_ = pv118_2_;
  assign pv151_3_ = new_n_n63_;
  assign pv183_11_ = new_n_n33_;
  assign pv199_7_ = new_n_n24_;
  assign new_n_n190_ = pv16_6_;
  assign new_n_n178_ = pv16_15_;
  assign new_n_n161_ = pv40_10_;
  assign new_n_n153_ = pv52_15_;
  assign new_n_n102_ = pv88_5_;
  assign new_n_n108_ = pv88_14_;
  assign new_n_n104_ = pv100_15_;
  assign new_n_n89_ = pv118_1_;
  assign new_n_n68_ = pv128_0_;
  assign pv151_2_ = new_n_n64_;
  assign pv167_10_ = new_n_n46_;
  assign pv183_12_ = new_n_n9_;
  assign pv199_6_ = new_n_n25_;
  assign new_n_n200_ = pv4_0_;
  assign new_n_n162_ = pv52_9_;
  assign new_n_n111_ = pv88_11_;
  assign new_n_n120_ = pv100_3_;
  assign new_n_n112_ = pv100_10_;
  assign new_n_n83_ = pv121_2_;
  assign new_n_n75_ = pv132_0_;
  assign pv167_4_ = new_n_n14_;
  assign pv199_1_ = new_n_n29_;
  assign new_n_n198_ = pv4_1_;
  assign new_n_n186_ = pv28_9_;
  assign new_n_n128_ = pv64_1_;
  assign new_n_n81_ = pv121_3_;
  assign pv167_5_ = new_n_n50_;
  assign pv199_0_ = new_n_n2_;
  assign new_n_n185_ = pv16_10_;
  assign new_n_n189_ = pv28_6_;
  assign new_n_n119_ = pv100_5_;
  assign pv167_2_ = new_n_n52_;
  assign pv199_3_ = new_n_n27_;
  assign new_n_n183_ = pv16_11_;
  assign new_n_n187_ = pv28_7_;
  assign new_n_n113_ = pv88_10_;
  assign new_n_n117_ = pv100_6_;
  assign new_n_n110_ = pv100_11_;
  assign new_n_n76_ = pv121_1_;
  assign pv167_3_ = new_n_n51_;
  assign pv199_2_ = new_n_n28_;
  assign new_n_n131_ = pv76_14_;
  assign pv167_8_ = new_n_n13_;
  assign pv199_14_ = new_n_n19_;
  assign new_n_n191_ = pv28_5_;
  assign new_n_n127_ = pv64_5_;
  assign new_n_n129_ = pv76_15_;
  assign pv167_9_ = new_n_n47_;
  assign pv199_15_ = new_n_n18_;
  assign new_n_n194_ = pv28_2_;
  assign new_n_n147_ = pv64_2_;
  assign new_n_n124_ = pv100_1_;
  assign pv167_6_ = new_n_n49_;
  assign pv199_12_ = new_n_n6_;
  assign new_n_n192_ = pv28_3_;
  assign new_n_n145_ = pv64_3_;
  assign new_n_n122_ = pv100_2_;
  assign pv167_7_ = new_n_n48_;
  assign pv199_13_ = new_n_n20_;
  assign new_n_n172_ = pv52_1_;
  assign new_n_n136_ = pv76_10_;
  assign new_n_n98_ = pv103_2_;
  assign new_n_n84_ = pv124_1_;
  assign pv199_10_ = new_n_n22_;
  assign new_n_n196_ = pv28_1_;
  assign new_n_n126_ = pv64_9_;
  assign new_n_n134_ = pv76_11_;
  assign new_n_n96_ = pv103_3_;
  assign new_n_n82_ = pv124_2_;
  assign pv199_11_ = new_n_n21_;
  assign new_n_n168_ = pv52_3_;
  assign new_n_n142_ = pv64_6_;
  assign new_n_n130_ = pv64_15_;
  assign new_n_n170_ = pv52_2_;
  assign new_n_n140_ = pv64_7_;
  assign new_n_n133_ = pv76_13_;
  assign new_n_n167_ = pv52_5_;
  assign new_n_n115_ = pv100_7_;
  assign new_n_n92_ = pv112_2_;
  assign pv167_0_ = new_n_n4_;
  assign pv183_6_ = new_n_n37_;
  assign new_n_n94_ = pv112_1_;
  assign new_n_n69_ = pv132_3_;
  assign new_n_n105_ = pv133_0_;
  assign pv167_1_ = new_n_n53_;
  assign pv183_7_ = new_n_n36_;
  assign new_n_n163_ = pv52_7_;
  assign new_n_n114_ = pv100_9_;
  assign new_n_n71_ = pv132_2_;
  assign pv183_8_ = new_n_n10_;
  assign new_n_n152_ = pv40_1_;
  assign new_n_n165_ = pv52_6_;
  assign new_n_n79_ = pv103_1_;
  assign new_n_n90_ = pv112_3_;
  assign new_n_n73_ = pv132_1_;
  assign pv183_9_ = new_n_n35_;
  assign new_n_n176_ = pv16_1_;
  assign new_n_n171_ = pv40_2_;
  assign new_n_n139_ = pv76_7_;
  assign new_n_n99_ = pv106_1_;
  assign pv151_5_ = new_n_n62_;
  assign pv151_14_ = new_n_n55_;
  assign pv183_2_ = new_n_n40_;
  assign pv183_13_ = new_n_n32_;
  assign new_n_n169_ = pv40_3_;
  assign new_n_n137_ = pv64_10_;
  assign new_n_n141_ = pv76_6_;
  assign new_n_n97_ = pv106_2_;
  assign pv151_4_ = new_n_n17_;
  assign pv151_15_ = new_n_n54_;
  assign pv183_3_ = new_n_n39_;
  assign pv183_14_ = new_n_n31_;
  assign new_n_n193_ = pv16_3_;
  assign new_n_n177_ = pv28_15_;
  assign new_n_n143_ = pv76_5_;
  assign new_n_n95_ = pv106_3_;
  assign pv151_7_ = new_n_n60_;
  assign pv151_12_ = new_n_n15_;
  assign pv183_4_ = new_n_n11_;
  assign pv183_15_ = new_n_n30_;
  assign new_n_n195_ = pv16_2_;
  assign new_n_n151_ = pv40_5_;
  assign new_n_n103_ = pv88_1_;
  assign pv151_6_ = new_n_n61_;
  assign pv151_13_ = new_n_n56_;
  assign pv183_5_ = new_n_n38_;
  assign new_n_n181_ = pv28_13_;
  assign new_n_n166_ = pv40_6_;
  assign new_n_n125_ = pv64_13_;
  assign new_n_n77_ = pv115_1_;
  assign pv151_9_ = new_n_n59_;
  assign pv151_10_ = new_n_n58_;
  assign pv167_15_ = new_n_n42_;
  assign new_n_n179_ = pv28_14_;
  assign new_n_n164_ = pv40_7_;
  assign new_n_n132_ = pv64_14_;
  assign pv151_8_ = new_n_n16_;
  assign pv151_11_ = new_n_n57_;
  assign new_n_n182_ = pv28_11_;
  assign new_n_n135_ = pv64_11_;
  assign new_n_n138_ = pv76_9_;
  assign new_n_n86_ = pv115_3_;
  assign new_n_n80_ = pv124_3_;
  assign pv135_1_ = new_n_n66_;
  assign pv183_0_ = new_n_n3_;
  assign new_n_n150_ = pv40_9_;
  assign new_n_n88_ = pv115_2_;
  assign pv135_0_ = new_n_n67_;
  assign pv183_1_ = new_n_n41_;
  assign new_n_n55_ = new_nv224_ | new_n_n180_ | new_nv225_;
  assign new_nv236_ = new_n_n164_ & new_n_n165_;
  assign new_nv247_ = new_n_n3_ & new_n_n157_ & new_n_n153_ & new_n_n155_;
  assign new_n_n46_ = new_nv242_ | new_n_n161_ | new_nv243_;
  assign new_nv257_ = new_n_n142_ & new_n_n143_;
  assign new_nv268_ = new_n_n134_ & new_n_n9_;
  assign new_n_n54_ = new_nv226_ | new_n_n178_;
  assign new_nv235_ = new_n_n13_ & new_n_n167_ & new_n_n163_ & new_n_n165_;
  assign new_nv248_ = new_n_n154_ & new_n_n155_;
  assign new_n_n47_ = new_nv241_ | new_n_n150_ | new_nv239_ | new_nv240_;
  assign new_nv258_ = new_n_n141_ & new_n_n140_ & new_n_n143_;
  assign new_nv267_ = new_n_n9_ & new_n_n136_ & new_n_n134_;
  assign new_nv217_ = new_n_n15_ & new_n_n186_ & new_n_n182_ & new_n_n184_;
  assign new_n_n64_ = new_nv206_ | new_n_n195_ | new_nv207_;
  assign new_nv249_ = new_n_n3_ & new_n_n155_ & new_n_n153_;
  assign new_n_n44_ = new_nv247_ | new_n_n149_ | new_nv245_ | new_nv246_;
  assign new_nv255_ = new_n_n11_ & new_n_n146_ & new_n_n144_;
  assign new_nv266_ = new_n_n135_ & new_n_n136_;
  assign new_nv218_ = new_n_n183_ & new_n_n184_;
  assign new_n_n65_ = new_nv205_ | new_n_n176_ | new_nv203_ | new_nv204_;
  assign new_nv250_ = new_n_n153_ & new_n_n3_;
  assign new_n_n45_ = new_nv244_ | new_n_n159_;
  assign new_nv256_ = new_n_n144_ & new_n_n11_;
  assign new_nv265_ = new_n_n9_ & new_n_n138_ & new_n_n134_ & new_n_n136_;
  assign new_nv208_ = new_n_n192_ & new_n_n17_;
  assign new_n_n53_ = new_nv229_ | new_n_n152_ | new_nv227_ | new_nv228_;
  assign new_n_n42_ = new_nv250_ | new_n_n154_;
  assign new_nv261_ = new_n_n10_ & new_n_n141_ & new_n_n139_;
  assign new_nv272_ = new_n_n130_ & new_n_n131_;
  assign new_nv327_ = new_n_n72_ & new_n_n73_;
  assign new_nv200_ = new_n_n199_ & new_n_n200_;
  assign new_nv207_ = new_n_n17_ & new_n_n194_ & new_n_n192_;
  assign new_n_n52_ = new_nv230_ | new_n_n171_ | new_nv231_;
  assign new_n_n43_ = new_nv248_ | new_n_n156_ | new_nv249_;
  assign new_nv262_ = new_n_n139_ & new_n_n10_;
  assign new_nv271_ = new_n_n2_ & new_n_n133_ & new_n_n129_ & new_n_n131_;
  assign new_n_n51_ = new_nv232_ | new_n_n169_;
  assign new_nv252_ = new_n_n146_ & new_n_n145_ & new_n_n148_;
  assign new_nv259_ = new_n_n10_ & new_n_n143_ & new_n_n139_ & new_n_n141_;
  assign new_nv270_ = new_n_n131_ & new_n_n130_ & new_n_n133_;
  assign new_n_n50_ = new_nv235_ | new_n_n151_ | new_nv233_ | new_nv234_;
  assign new_nv251_ = new_n_n147_ & new_n_n148_;
  assign new_nv260_ = new_n_n140_ & new_n_n141_;
  assign new_nv269_ = new_n_n132_ & new_n_n133_;
  assign new_n_n67_ = new_nv200_ | new_n_n197_ | new_nv201_;
  assign new_nv212_ = new_n_n188_ & new_n_n189_;
  assign new_nv223_ = new_n_n4_ & new_n_n181_ & new_n_n177_ & new_n_n179_;
  assign new_n_n58_ = new_nv218_ | new_n_n185_ | new_nv219_;
  assign new_nv233_ = new_n_n166_ & new_n_n167_;
  assign new_nv244_ = new_n_n158_ & new_n_n12_;
  assign new_nv331_ = new_n_n105_ & new_n_n71_ & new_n_n69_;
  assign new_n_n66_ = new_nv202_ | new_n_n199_;
  assign new_nv211_ = new_n_n16_ & new_n_n191_ & new_n_n187_ & new_n_n189_;
  assign new_nv224_ = new_n_n178_ & new_n_n179_;
  assign new_n_n59_ = new_nv217_ | new_n_n174_ | new_nv215_ | new_nv216_;
  assign new_nv234_ = new_n_n165_ & new_n_n164_ & new_n_n167_;
  assign new_nv243_ = new_n_n12_ & new_n_n160_ & new_n_n158_;
  assign new_nv330_ = new_n_n70_ & new_n_n71_;
  assign new_nv201_ = new_n_n5_ & new_n_n200_ & new_n_n198_;
  assign new_nv210_ = new_n_n189_ & new_n_n188_ & new_n_n191_;
  assign new_nv225_ = new_n_n4_ & new_n_n179_ & new_n_n177_;
  assign new_n_n56_ = new_nv223_ | new_n_n173_ | new_nv221_ | new_nv222_;
  assign new_nv231_ = new_n_n14_ & new_n_n170_ & new_n_n168_;
  assign new_nv242_ = new_n_n159_ & new_n_n160_;
  assign new_nv329_ = new_n_n105_ & new_n_n73_ & new_n_n69_ & new_n_n71_;
  assign new_nv202_ = new_n_n198_ & new_n_n5_;
  assign new_nv209_ = new_n_n190_ & new_n_n191_;
  assign new_nv226_ = new_n_n177_ & new_n_n4_;
  assign new_n_n57_ = new_nv220_ | new_n_n183_;
  assign new_nv232_ = new_n_n168_ & new_n_n14_;
  assign new_nv241_ = new_n_n12_ & new_n_n162_ & new_n_n158_ & new_n_n160_;
  assign new_nv328_ = new_n_n71_ & new_n_n70_ & new_n_n73_;
  assign new_nv205_ = new_n_n17_ & new_n_n196_ & new_n_n192_ & new_n_n194_;
  assign new_nv216_ = new_n_n184_ & new_n_n183_ & new_n_n186_;
  assign new_nv219_ = new_n_n15_ & new_n_n184_ & new_n_n182_;
  assign new_n_n62_ = new_nv211_ | new_n_n175_ | new_nv209_ | new_nv210_;
  assign new_nv229_ = new_n_n14_ & new_n_n172_ & new_n_n168_ & new_n_n170_;
  assign new_nv240_ = new_n_n160_ & new_n_n159_ & new_n_n162_;
  assign new_nv253_ = new_n_n11_ & new_n_n148_ & new_n_n144_ & new_n_n146_;
  assign new_nv264_ = new_n_n136_ & new_n_n135_ & new_n_n138_;
  assign new_n_n3_ = new_nv330_ | new_n_n72_ | new_nv331_;
  assign new_nv206_ = new_n_n193_ & new_n_n194_;
  assign new_nv215_ = new_n_n185_ & new_n_n186_;
  assign new_nv220_ = new_n_n182_ & new_n_n15_;
  assign new_n_n63_ = new_nv208_ | new_n_n193_;
  assign new_nv230_ = new_n_n169_ & new_n_n170_;
  assign new_nv239_ = new_n_n161_ & new_n_n162_;
  assign new_nv254_ = new_n_n145_ & new_n_n146_;
  assign new_nv263_ = new_n_n137_ & new_n_n138_;
  assign new_n_n4_ = new_nv329_ | new_n_n74_ | new_nv327_ | new_nv328_;
  assign new_nv203_ = new_n_n195_ & new_n_n196_;
  assign new_nv214_ = new_n_n187_ & new_n_n16_;
  assign new_nv221_ = new_n_n180_ & new_n_n181_;
  assign new_n_n60_ = new_nv214_ | new_n_n188_;
  assign new_nv227_ = new_n_n171_ & new_n_n172_;
  assign new_nv238_ = new_n_n163_ & new_n_n13_;
  assign new_nv245_ = new_n_n156_ & new_n_n157_;
  assign new_n_n48_ = new_nv238_ | new_n_n164_;
  assign new_n_n5_ = new_nv323_ | new_nv324_ | new_nv326_ | new_n_n68_ | new_nv325_;
  assign new_nv204_ = new_n_n194_ & new_n_n193_ & new_n_n196_;
  assign new_nv213_ = new_n_n16_ & new_n_n189_ & new_n_n187_;
  assign new_nv222_ = new_n_n179_ & new_n_n178_ & new_n_n181_;
  assign new_n_n61_ = new_nv212_ | new_n_n190_ | new_nv213_;
  assign new_nv228_ = new_n_n170_ & new_n_n169_ & new_n_n172_;
  assign new_nv237_ = new_n_n13_ & new_n_n165_ & new_n_n163_;
  assign new_nv246_ = new_n_n155_ & new_n_n154_ & new_n_n157_;
  assign new_n_n49_ = new_nv236_ | new_n_n166_ | new_nv237_;
  assign new_nv332_ = new_n_n69_ & new_n_n105_;
  assign new_n_n38_ = new_nv259_ | new_n_n127_ | new_nv257_ | new_nv258_;
  assign new_nv277_ = new_n_n8_ & new_n_n124_ & new_n_n120_ & new_n_n122_;
  assign new_nv288_ = new_n_n112_ & new_n_n111_ & new_n_n114_;
  assign new_n_n29_ = new_nv277_ | new_n_n103_ | new_nv275_ | new_nv276_;
  assign new_n_n18_ = new_nv298_ | new_n_n106_;
  assign new_n_n39_ = new_nv256_ | new_n_n145_;
  assign new_nv278_ = new_n_n121_ & new_n_n122_;
  assign new_nv287_ = new_n_n113_ & new_n_n114_;
  assign new_n_n28_ = new_nv278_ | new_n_n123_ | new_nv279_;
  assign new_n_n19_ = new_nv296_ | new_n_n108_ | new_nv297_;
  assign new_n_n40_ = new_nv254_ | new_n_n147_ | new_nv255_;
  assign new_nv279_ = new_n_n8_ & new_n_n122_ & new_n_n120_;
  assign new_nv290_ = new_n_n111_ & new_n_n112_;
  assign new_nv297_ = new_n_n105_ & new_n_n107_ & new_n_n104_;
  assign new_n_n20_ = new_nv295_ | new_n_n100_ | new_nv293_ | new_nv294_;
  assign new_n_n41_ = new_nv253_ | new_n_n128_ | new_nv251_ | new_nv252_;
  assign new_nv280_ = new_n_n120_ & new_n_n8_;
  assign new_nv289_ = new_n_n6_ & new_n_n114_ & new_n_n110_ & new_n_n112_;
  assign new_nv298_ = new_n_n104_ & new_n_n105_;
  assign new_n_n21_ = new_nv292_ | new_n_n111_;
  assign new_n_n2_ = new_nv332_ | new_n_n70_;
  assign new_nv274_ = new_n_n129_ & new_n_n2_;
  assign new_nv305_ = new_n_n93_ & new_n_n94_;
  assign new_nv316_ = new_n_n85_ & new_n_n2_;
  assign new_n_n13_ = new_nv308_ | new_n_n93_ | new_nv309_;
  assign new_nv326_ = new_n_n105_ & new_n_n75_ & new_n_n71_ & new_n_n73_ & new_n_n69_;
  assign new_nv273_ = new_n_n2_ & new_n_n131_ & new_n_n129_;
  assign new_nv306_ = new_n_n92_ & new_n_n91_ & new_n_n94_;
  assign new_nv315_ = new_n_n2_ & new_n_n87_ & new_n_n85_;
  assign new_n_n12_ = new_nv310_ | new_n_n91_;
  assign new_nv325_ = new_n_n71_ & new_n_n70_ & new_n_n73_ & new_n_n75_;
  assign new_nv307_ = new_n_n3_ & new_n_n94_ & new_n_n90_ & new_n_n92_;
  assign new_nv318_ = new_n_n82_ & new_n_n81_ & new_n_n84_;
  assign new_n_n15_ = new_nv304_ | new_n_n96_;
  assign new_nv324_ = new_n_n73_ & new_n_n72_ & new_n_n75_;
  assign new_nv308_ = new_n_n91_ & new_n_n92_;
  assign new_nv317_ = new_n_n83_ & new_n_n84_;
  assign new_n_n14_ = new_nv307_ | new_n_n78_ | new_nv305_ | new_nv306_;
  assign new_nv323_ = new_n_n74_ & new_n_n75_;
  assign new_nv291_ = new_n_n6_ & new_n_n112_ & new_n_n110_;
  assign new_n_n26_ = new_nv283_ | new_n_n102_ | new_nv281_ | new_nv282_;
  assign new_nv301_ = new_n_n4_ & new_n_n99_ & new_n_n95_ & new_n_n97_;
  assign new_nv312_ = new_n_n87_ & new_n_n86_ & new_n_n89_;
  assign new_n_n17_ = new_nv301_ | new_n_n79_ | new_nv299_ | new_nv300_;
  assign new_n_n6_ = new_nv322_ | new_n_n81_;
  assign new_nv292_ = new_n_n110_ & new_n_n6_;
  assign new_n_n27_ = new_nv280_ | new_n_n121_;
  assign new_nv302_ = new_n_n96_ & new_n_n97_;
  assign new_nv311_ = new_n_n88_ & new_n_n89_;
  assign new_n_n16_ = new_nv302_ | new_n_n98_ | new_nv303_;
  assign new_n_n7_ = new_nv320_ | new_n_n83_ | new_nv321_;
  assign new_n_n33_ = new_nv268_ | new_n_n135_;
  assign new_nv282_ = new_n_n117_ & new_n_n116_ & new_n_n119_;
  assign new_nv303_ = new_n_n4_ & new_n_n97_ & new_n_n95_;
  assign new_nv314_ = new_n_n86_ & new_n_n87_;
  assign new_nv321_ = new_n_n105_ & new_n_n82_ & new_n_n80_;
  assign new_n_n8_ = new_nv319_ | new_n_n76_ | new_nv317_ | new_nv318_;
  assign new_n_n32_ = new_nv271_ | new_n_n125_ | new_nv269_ | new_nv270_;
  assign new_nv281_ = new_n_n118_ & new_n_n119_;
  assign new_nv304_ = new_n_n95_ & new_n_n4_;
  assign new_nv313_ = new_n_n2_ & new_n_n89_ & new_n_n85_ & new_n_n87_;
  assign new_nv322_ = new_n_n80_ & new_n_n105_;
  assign new_n_n9_ = new_nv316_ | new_n_n86_;
  assign new_n_n34_ = new_nv266_ | new_n_n137_ | new_nv267_;
  assign new_n_n31_ = new_nv272_ | new_n_n132_ | new_nv273_;
  assign new_nv284_ = new_n_n116_ & new_n_n117_;
  assign new_nv295_ = new_n_n105_ & new_n_n109_ & new_n_n104_ & new_n_n107_;
  assign new_n_n22_ = new_nv290_ | new_n_n113_ | new_nv291_;
  assign new_nv319_ = new_n_n105_ & new_n_n84_ & new_n_n80_ & new_n_n82_;
  assign new_n_n10_ = new_nv314_ | new_n_n88_ | new_nv315_;
  assign new_n_n35_ = new_nv265_ | new_n_n126_ | new_nv263_ | new_nv264_;
  assign new_n_n30_ = new_nv274_ | new_n_n130_;
  assign new_nv283_ = new_n_n7_ & new_n_n119_ & new_n_n115_ & new_n_n117_;
  assign new_nv296_ = new_n_n106_ & new_n_n107_;
  assign new_n_n23_ = new_nv289_ | new_n_n101_ | new_nv287_ | new_nv288_;
  assign new_nv320_ = new_n_n81_ & new_n_n82_;
  assign new_n_n11_ = new_nv313_ | new_n_n77_ | new_nv311_ | new_nv312_;
  assign new_n_n36_ = new_nv262_ | new_n_n140_;
  assign new_nv275_ = new_n_n123_ & new_n_n124_;
  assign new_nv286_ = new_n_n115_ & new_n_n7_;
  assign new_nv293_ = new_n_n108_ & new_n_n109_;
  assign new_n_n24_ = new_nv286_ | new_n_n116_;
  assign new_nv299_ = new_n_n98_ & new_n_n99_;
  assign new_nv310_ = new_n_n90_ & new_n_n3_;
  assign new_n_n37_ = new_nv260_ | new_n_n142_ | new_nv261_;
  assign new_nv276_ = new_n_n122_ & new_n_n121_ & new_n_n124_;
  assign new_nv285_ = new_n_n7_ & new_n_n117_ & new_n_n115_;
  assign new_nv294_ = new_n_n107_ & new_n_n106_ & new_n_n109_;
  assign new_n_n25_ = new_nv284_ | new_n_n118_ | new_nv285_;
  assign new_nv300_ = new_n_n97_ & new_n_n96_ & new_n_n99_;
  assign new_nv309_ = new_n_n3_ & new_n_n92_ & new_n_n90_;
endmodule


