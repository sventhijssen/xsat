// Benchmark "top" written by ABC on Fri Mar 31 12:10:02 2023

module top ( 
    pv144_18_, pv126_20_, pv126_31_, pv94_30_, pv126_9_, pv129_0_,
    pv94_31_, pv144_19_, pv94_10_, pv94_21_, pv126_7_, pv126_10_,
    pv144_27_, pv176_31_, pv190_0_, pv94_11_, pv94_20_, pv126_8_,
    pv144_28_, pv176_30_, pv30_18_, pv30_29_, pv126_5_, pv144_29_,
    pv30_19_, pv30_28_, pv126_6_, pv128_0_, pv190_1_, pv30_9_, pv62_2_,
    pv64_0_, pv126_14_, pv126_27_, pv176_8_, pv176_22_, pv188_23_, pv30_8_,
    pv62_3_, pv126_13_, pv126_28_, pv176_7_, pv176_23_, pv178_1_,
    pv188_24_, pv30_7_, pv62_0_, pv126_12_, pv126_25_, pv176_6_, pv176_20_,
    pv178_0_, pv188_25_, pv30_6_, pv62_1_, pv63_0_, pv126_11_, pv126_26_,
    pv176_5_, pv176_21_, pv188_26_, pv30_5_, pv62_6_, pv94_7_, pv126_18_,
    pv126_23_, pv176_13_, pv188_27_, pv30_4_, pv62_7_, pv94_6_, pv126_17_,
    pv126_24_, pv176_12_, pv188_28_, pv30_3_, pv62_4_, pv94_9_, pv126_16_,
    pv126_21_, pv126_30_, pv130_0_, pv176_11_, pv188_29_, pv30_2_, pv62_5_,
    pv94_8_, pv126_15_, pv126_22_, pv176_9_, pv176_10_, pv30_30_, pv62_15_,
    pv62_26_, pv94_3_, pv176_0_, pv176_17_, pv30_31_, pv62_16_, pv62_25_,
    pv94_2_, pv176_16_, pv201_0_, pv62_8_, pv62_17_, pv62_28_, pv94_5_,
    pv176_15_, pv176_28_, pv201_1_, pv62_9_, pv62_18_, pv62_27_, pv94_4_,
    pv126_19_, pv176_14_, pv176_29_, pv191_31_, pv201_2_, pv62_19_,
    pv176_4_, pv176_26_, pv62_29_, pv176_3_, pv176_27_, pv188_31_,
    pv126_29_, pv176_2_, pv176_19_, pv176_24_, pv188_30_, pv176_1_,
    pv176_18_, pv176_25_, pv188_22_, pv30_16_, pv30_27_, pv94_14_,
    pv94_25_, pv126_3_, pv127_0_, pv144_23_, pv201_7_, pv30_17_, pv30_26_,
    pv62_30_, pv94_15_, pv94_24_, pv126_4_, pv144_24_, pv30_14_, pv30_25_,
    pv62_20_, pv94_12_, pv94_23_, pv126_1_, pv144_25_, pv30_15_, pv30_24_,
    pv62_10_, pv94_13_, pv94_22_, pv126_2_, pv144_26_, pv30_12_, pv30_23_,
    pv62_11_, pv62_22_, pv94_18_, pv94_29_, pv201_3_, pv30_13_, pv30_22_,
    pv62_12_, pv62_21_, pv94_19_, pv94_28_, pv126_0_, pv144_20_, pv144_31_,
    pv201_4_, pv30_10_, pv30_21_, pv62_13_, pv62_24_, pv62_31_, pv94_16_,
    pv94_27_, pv144_21_, pv144_30_, pv193_1_, pv201_5_, pv30_11_, pv30_20_,
    pv62_14_, pv62_23_, pv94_17_, pv94_26_, pv144_22_, pv193_0_, pv201_6_,
    pv202_0_  );
  input  pv144_18_, pv126_20_, pv126_31_, pv94_30_, pv126_9_, pv129_0_,
    pv94_31_, pv144_19_, pv94_10_, pv94_21_, pv126_7_, pv126_10_,
    pv144_27_, pv176_31_, pv190_0_, pv94_11_, pv94_20_, pv126_8_,
    pv144_28_, pv176_30_, pv30_18_, pv30_29_, pv126_5_, pv144_29_,
    pv30_19_, pv30_28_, pv126_6_, pv128_0_, pv190_1_, pv30_9_, pv62_2_,
    pv64_0_, pv126_14_, pv126_27_, pv176_8_, pv176_22_, pv188_23_, pv30_8_,
    pv62_3_, pv126_13_, pv126_28_, pv176_7_, pv176_23_, pv178_1_,
    pv188_24_, pv30_7_, pv62_0_, pv126_12_, pv126_25_, pv176_6_, pv176_20_,
    pv178_0_, pv188_25_, pv30_6_, pv62_1_, pv63_0_, pv126_11_, pv126_26_,
    pv176_5_, pv176_21_, pv188_26_, pv30_5_, pv62_6_, pv94_7_, pv126_18_,
    pv126_23_, pv176_13_, pv188_27_, pv30_4_, pv62_7_, pv94_6_, pv126_17_,
    pv126_24_, pv176_12_, pv188_28_, pv30_3_, pv62_4_, pv94_9_, pv126_16_,
    pv126_21_, pv126_30_, pv130_0_, pv176_11_, pv188_29_, pv30_2_, pv62_5_,
    pv94_8_, pv126_15_, pv126_22_, pv176_9_, pv176_10_, pv30_30_, pv62_15_,
    pv62_26_, pv94_3_, pv176_0_, pv176_17_, pv30_31_, pv62_16_, pv62_25_,
    pv94_2_, pv176_16_, pv201_0_, pv62_8_, pv62_17_, pv62_28_, pv94_5_,
    pv176_15_, pv176_28_, pv201_1_, pv62_9_, pv62_18_, pv62_27_, pv94_4_,
    pv126_19_, pv176_14_, pv176_29_, pv191_31_, pv201_2_, pv62_19_,
    pv176_4_, pv176_26_, pv62_29_, pv176_3_, pv176_27_, pv188_31_,
    pv126_29_, pv176_2_, pv176_19_, pv176_24_, pv188_30_, pv176_1_,
    pv176_18_, pv176_25_, pv188_22_, pv30_16_, pv30_27_, pv94_14_,
    pv94_25_, pv126_3_, pv127_0_, pv144_23_, pv201_7_, pv30_17_, pv30_26_,
    pv62_30_, pv94_15_, pv94_24_, pv126_4_, pv144_24_, pv30_14_, pv30_25_,
    pv62_20_, pv94_12_, pv94_23_, pv126_1_, pv144_25_, pv30_15_, pv30_24_,
    pv62_10_, pv94_13_, pv94_22_, pv126_2_, pv144_26_, pv30_12_, pv30_23_,
    pv62_11_, pv62_22_, pv94_18_, pv94_29_, pv201_3_, pv30_13_, pv30_22_,
    pv62_12_, pv62_21_, pv94_19_, pv94_28_, pv126_0_, pv144_20_, pv144_31_,
    pv201_4_, pv30_10_, pv30_21_, pv62_13_, pv62_24_, pv62_31_, pv94_16_,
    pv94_27_, pv144_21_, pv144_30_, pv193_1_, pv201_5_, pv30_11_, pv30_20_,
    pv62_14_, pv62_23_, pv94_17_, pv94_26_, pv144_22_, pv193_0_, pv201_6_;
  output pv202_0_;
  wire new_n_n73_, new_n_n92_, new_n_n116_, new_n_n119_, new_n_n105_,
    new_n_n84_, new_n_n148_, new_n_n74_, new_n_n129_, new_n_n143_,
    new_n_n104_, new_n_n97_, new_n_n78_, new_n_n48_, new_n_n20_,
    new_n_n138_, new_n_n124_, new_n_n98_, new_n_n68_, new_n_n35_,
    new_n_n189_, new_n_n211_, new_n_n103_, new_n_n79_, new_n_n206_,
    new_n_n184_, new_n_n99_, new_n_n117_, new_n_n23_, new_n_n201_,
    new_n_n165_, new_n_n181_, new_n_n95_, new_n_n114_, new_n_n54_,
    new_n_n39_, new_n_n30_, new_n_n194_, new_n_n166_, new_n_n107_,
    new_n_n88_, new_n_n60_, new_n_n44_, new_n_n49_, new_n_n28_,
    new_n_n200_, new_n_n182_, new_n_n96_, new_n_n113_, new_n_n55_,
    new_n_n40_, new_n_n34_, new_n_n31_, new_n_n195_, new_n_n213_,
    new_n_n150_, new_n_n106_, new_n_n89_, new_n_n59_, new_n_n43_,
    new_n_n25_, new_n_n199_, new_n_n163_, new_n_n136_, new_n_n93_,
    new_n_n112_, new_n_n63_, new_n_n26_, new_n_n196_, new_n_n168_,
    new_n_n131_, new_n_n109_, new_n_n90_, new_n_n52_, new_n_n24_,
    new_n_n198_, new_n_n164_, new_n_n137_, new_n_n94_, new_n_n111_,
    new_n_n87_, new_n_n82_, new_n_n62_, new_n_n27_, new_n_n197_,
    new_n_n167_, new_n_n130_, new_n_n108_, new_n_n91_, new_n_n61_,
    new_n_n53_, new_n_n183_, new_n_n172_, new_n_n153_, new_n_n134_,
    new_n_n66_, new_n_n65_, new_n_n212_, new_n_n158_, new_n_n177_,
    new_n_n133_, new_n_n50_, new_n_n85_, new_n_n162_, new_n_n173_,
    new_n_n152_, new_n_n135_, new_n_n64_, new_n_n36_, new_n_n83_,
    new_n_n169_, new_n_n157_, new_n_n178_, new_n_n132_, new_n_n110_,
    new_n_n51_, new_n_n47_, new_n_n16_, new_n_n32_, new_n_n174_,
    new_n_n56_, new_n_n37_, new_n_n179_, new_n_n58_, new_n_n46_,
    new_n_n22_, new_n_n115_, new_n_n57_, new_n_n42_, new_n_n38_,
    new_n_n21_, new_n_n81_, new_n_n41_, new_n_n45_, new_n_n29_,
    new_n_n190_, new_n_n210_, new_n_n127_, new_n_n145_, new_n_n102_,
    new_n_n86_, new_n_n76_, new_n_n17_, new_n_n205_, new_n_n185_,
    new_n_n151_, new_n_n140_, new_n_n122_, new_n_n100_, new_n_n70_,
    new_n_n191_, new_n_n209_, new_n_n156_, new_n_n128_, new_n_n144_,
    new_n_n149_, new_n_n77_, new_n_n204_, new_n_n186_, new_n_n161_,
    new_n_n139_, new_n_n123_, new_n_n101_, new_n_n69_, new_n_n192_,
    new_n_n208_, new_n_n170_, new_n_n155_, new_n_n125_, new_n_n147_,
    new_n_n33_, new_n_n203_, new_n_n187_, new_n_n160_, new_n_n175_,
    new_n_n142_, new_n_n120_, new_n_n118_, new_n_n72_, new_n_n80_,
    new_n_n18_, new_n_n193_, new_n_n207_, new_n_n171_, new_n_n154_,
    new_n_n180_, new_n_n126_, new_n_n146_, new_n_n75_, new_n_n67_,
    new_n_n13_, new_n_n19_, new_n_n202_, new_n_n188_, new_n_n159_,
    new_n_n176_, new_n_n141_, new_n_n121_, new_n_n71_, new_n_n14_,
    new_n_n15_, new_nv230_, new_nv234_, new_nv233_, new_nv232_, new_nv231_,
    new_n_n12_, new_nv237_, new_nv236_, new_nv235_, new_nv207_, new_n_n8_,
    new_nv218_, new_nv229_, new_n_n9_, new_nv219_, new_nv228_, new_nv209_,
    new_n_n5_, new_nv227_, new_nv208_, new_nv217_, new_nv226_, new_n_n7_,
    new_n_n2_, new_n_n6_, new_n_n3_, new_n_n10_, new_nv212_, new_n_n4_,
    new_n_n11_, new_nv213_, new_nv222_, new_nv210_, new_nv221_, new_nv211_,
    new_nv220_;
  assign new_n_n73_ = pv144_18_;
  assign new_n_n92_ = pv126_20_;
  assign new_n_n116_ = pv126_31_;
  assign new_n_n119_ = pv94_30_;
  assign new_n_n105_ = pv126_9_;
  assign new_n_n84_ = pv129_0_;
  assign new_n_n148_ = pv94_31_;
  assign new_n_n74_ = pv144_19_;
  assign new_n_n129_ = pv94_10_;
  assign new_n_n143_ = pv94_21_;
  assign new_n_n104_ = pv126_7_;
  assign new_n_n97_ = pv126_10_;
  assign new_n_n78_ = pv144_27_;
  assign new_n_n48_ = pv176_31_;
  assign new_n_n20_ = pv190_0_;
  assign new_n_n138_ = pv94_11_;
  assign new_n_n124_ = pv94_20_;
  assign new_n_n98_ = pv126_8_;
  assign new_n_n68_ = pv144_28_;
  assign new_n_n35_ = pv176_30_;
  assign new_n_n189_ = pv30_18_;
  assign new_n_n211_ = pv30_29_;
  assign new_n_n103_ = pv126_5_;
  assign new_n_n79_ = pv144_29_;
  assign new_n_n206_ = pv30_19_;
  assign new_n_n184_ = pv30_28_;
  assign new_n_n99_ = pv126_6_;
  assign new_n_n117_ = pv128_0_;
  assign new_n_n23_ = pv190_1_;
  assign new_n_n201_ = pv30_9_;
  assign new_n_n165_ = pv62_2_;
  assign new_n_n181_ = pv64_0_;
  assign new_n_n95_ = pv126_14_;
  assign new_n_n114_ = pv126_27_;
  assign new_n_n54_ = pv176_8_;
  assign new_n_n39_ = pv176_22_;
  assign new_n_n30_ = pv188_23_;
  assign new_n_n194_ = pv30_8_;
  assign new_n_n166_ = pv62_3_;
  assign new_n_n107_ = pv126_13_;
  assign new_n_n88_ = pv126_28_;
  assign new_n_n60_ = pv176_7_;
  assign new_n_n44_ = pv176_23_;
  assign new_n_n49_ = pv178_1_;
  assign new_n_n28_ = pv188_24_;
  assign new_n_n200_ = pv30_7_;
  assign new_n_n182_ = pv62_0_;
  assign new_n_n96_ = pv126_12_;
  assign new_n_n113_ = pv126_25_;
  assign new_n_n55_ = pv176_6_;
  assign new_n_n40_ = pv176_20_;
  assign new_n_n34_ = pv178_0_;
  assign new_n_n31_ = pv188_25_;
  assign new_n_n195_ = pv30_6_;
  assign new_n_n213_ = pv62_1_;
  assign new_n_n150_ = pv63_0_;
  assign new_n_n106_ = pv126_11_;
  assign new_n_n89_ = pv126_26_;
  assign new_n_n59_ = pv176_5_;
  assign new_n_n43_ = pv176_21_;
  assign new_n_n25_ = pv188_26_;
  assign new_n_n199_ = pv30_5_;
  assign new_n_n163_ = pv62_6_;
  assign new_n_n136_ = pv94_7_;
  assign new_n_n93_ = pv126_18_;
  assign new_n_n112_ = pv126_23_;
  assign new_n_n63_ = pv176_13_;
  assign new_n_n26_ = pv188_27_;
  assign new_n_n196_ = pv30_4_;
  assign new_n_n168_ = pv62_7_;
  assign new_n_n131_ = pv94_6_;
  assign new_n_n109_ = pv126_17_;
  assign new_n_n90_ = pv126_24_;
  assign new_n_n52_ = pv176_12_;
  assign new_n_n24_ = pv188_28_;
  assign new_n_n198_ = pv30_3_;
  assign new_n_n164_ = pv62_4_;
  assign new_n_n137_ = pv94_9_;
  assign new_n_n94_ = pv126_16_;
  assign new_n_n111_ = pv126_21_;
  assign new_n_n87_ = pv126_30_;
  assign new_n_n82_ = pv130_0_;
  assign new_n_n62_ = pv176_11_;
  assign new_n_n27_ = pv188_29_;
  assign new_n_n197_ = pv30_2_;
  assign new_n_n167_ = pv62_5_;
  assign new_n_n130_ = pv94_8_;
  assign new_n_n108_ = pv126_15_;
  assign new_n_n91_ = pv126_22_;
  assign new_n_n61_ = pv176_9_;
  assign new_n_n53_ = pv176_10_;
  assign new_n_n183_ = pv30_30_;
  assign new_n_n172_ = pv62_15_;
  assign new_n_n153_ = pv62_26_;
  assign new_n_n134_ = pv94_3_;
  assign new_n_n66_ = pv176_0_;
  assign new_n_n65_ = pv176_17_;
  assign new_n_n212_ = pv30_31_;
  assign new_n_n158_ = pv62_16_;
  assign new_n_n177_ = pv62_25_;
  assign new_n_n133_ = pv94_2_;
  assign new_n_n50_ = pv176_16_;
  assign new_n_n85_ = pv201_0_;
  assign new_n_n162_ = pv62_8_;
  assign new_n_n173_ = pv62_17_;
  assign new_n_n152_ = pv62_28_;
  assign new_n_n135_ = pv94_5_;
  assign new_n_n64_ = pv176_15_;
  assign new_n_n36_ = pv176_28_;
  assign new_n_n83_ = pv201_1_;
  assign new_n_n169_ = pv62_9_;
  assign new_n_n157_ = pv62_18_;
  assign new_n_n178_ = pv62_27_;
  assign new_n_n132_ = pv94_4_;
  assign new_n_n110_ = pv126_19_;
  assign new_n_n51_ = pv176_14_;
  assign new_n_n47_ = pv176_29_;
  assign new_n_n16_ = pv191_31_;
  assign new_n_n32_ = pv201_2_;
  assign new_n_n174_ = pv62_19_;
  assign new_n_n56_ = pv176_4_;
  assign new_n_n37_ = pv176_26_;
  assign new_n_n179_ = pv62_29_;
  assign new_n_n58_ = pv176_3_;
  assign new_n_n46_ = pv176_27_;
  assign new_n_n22_ = pv188_31_;
  assign new_n_n115_ = pv126_29_;
  assign new_n_n57_ = pv176_2_;
  assign new_n_n42_ = pv176_19_;
  assign new_n_n38_ = pv176_24_;
  assign new_n_n21_ = pv188_30_;
  assign new_n_n81_ = pv176_1_;
  assign new_n_n41_ = pv176_18_;
  assign new_n_n45_ = pv176_25_;
  assign new_n_n29_ = pv188_22_;
  assign new_n_n190_ = pv30_16_;
  assign new_n_n210_ = pv30_27_;
  assign new_n_n127_ = pv94_14_;
  assign new_n_n145_ = pv94_25_;
  assign new_n_n102_ = pv126_3_;
  assign new_n_n86_ = pv127_0_;
  assign new_n_n76_ = pv144_23_;
  assign new_n_n17_ = pv201_7_;
  assign new_n_n205_ = pv30_17_;
  assign new_n_n185_ = pv30_26_;
  assign new_n_n151_ = pv62_30_;
  assign new_n_n140_ = pv94_15_;
  assign new_n_n122_ = pv94_24_;
  assign new_n_n100_ = pv126_4_;
  assign new_n_n70_ = pv144_24_;
  assign new_n_n191_ = pv30_14_;
  assign new_n_n209_ = pv30_25_;
  assign new_n_n156_ = pv62_20_;
  assign new_n_n128_ = pv94_12_;
  assign new_n_n144_ = pv94_23_;
  assign new_n_n149_ = pv126_1_;
  assign new_n_n77_ = pv144_25_;
  assign new_n_n204_ = pv30_15_;
  assign new_n_n186_ = pv30_24_;
  assign new_n_n161_ = pv62_10_;
  assign new_n_n139_ = pv94_13_;
  assign new_n_n123_ = pv94_22_;
  assign new_n_n101_ = pv126_2_;
  assign new_n_n69_ = pv144_26_;
  assign new_n_n192_ = pv30_12_;
  assign new_n_n208_ = pv30_23_;
  assign new_n_n170_ = pv62_11_;
  assign new_n_n155_ = pv62_22_;
  assign new_n_n125_ = pv94_18_;
  assign new_n_n147_ = pv94_29_;
  assign new_n_n33_ = pv201_3_;
  assign pv202_0_ = new_n_n12_;
  assign new_n_n203_ = pv30_13_;
  assign new_n_n187_ = pv30_22_;
  assign new_n_n160_ = pv62_12_;
  assign new_n_n175_ = pv62_21_;
  assign new_n_n142_ = pv94_19_;
  assign new_n_n120_ = pv94_28_;
  assign new_n_n118_ = pv126_0_;
  assign new_n_n72_ = pv144_20_;
  assign new_n_n80_ = pv144_31_;
  assign new_n_n18_ = pv201_4_;
  assign new_n_n193_ = pv30_10_;
  assign new_n_n207_ = pv30_21_;
  assign new_n_n171_ = pv62_13_;
  assign new_n_n154_ = pv62_24_;
  assign new_n_n180_ = pv62_31_;
  assign new_n_n126_ = pv94_16_;
  assign new_n_n146_ = pv94_27_;
  assign new_n_n75_ = pv144_21_;
  assign new_n_n67_ = pv144_30_;
  assign new_n_n13_ = pv193_1_;
  assign new_n_n19_ = pv201_5_;
  assign new_n_n202_ = pv30_11_;
  assign new_n_n188_ = pv30_20_;
  assign new_n_n159_ = pv62_14_;
  assign new_n_n176_ = pv62_23_;
  assign new_n_n141_ = pv94_17_;
  assign new_n_n121_ = pv94_26_;
  assign new_n_n71_ = pv144_22_;
  assign new_n_n14_ = pv193_0_;
  assign new_n_n15_ = pv201_6_;
  assign new_nv230_ = new_nv229_ & new_n_n19_;
  assign new_nv234_ = new_nv233_ & new_n_n17_;
  assign new_nv233_ = new_n_n14_ & new_n_n15_;
  assign new_nv232_ = new_n_n17_ & new_n_n16_ & new_n_n15_;
  assign new_nv231_ = new_n_n2_ & new_n_n19_;
  assign new_n_n12_ = new_nv220_ | new_nv217_ | new_nv226_ | new_nv221_ | new_nv208_ | new_nv212_ | new_nv231_ | new_nv234_ | new_nv210_ | new_nv219_ | new_nv211_ | new_nv213_ | new_nv233_ | new_nv237_ | new_nv209_ | new_nv227_ | new_nv222_ | new_nv228_ | new_nv218_ | new_nv232_ | new_nv235_ | new_nv236_ | new_nv229_ | new_nv230_;
  assign new_nv237_ = new_n_n13_ & new_n_n17_;
  assign new_nv236_ = new_nv235_ & new_n_n17_;
  assign new_nv235_ = new_n_n13_ & new_n_n15_;
  assign new_nv207_ = ~new_n_n85_;
  assign new_n_n8_ = new_n_n91_ | new_n_n92_ | new_n_n93_ | new_n_n94_ | new_n_n97_ | new_n_n95_ | new_n_n96_ | new_n_n106_ | new_n_n117_ | new_n_n107_ | new_n_n101_ | new_n_n116_ | new_n_n100_ | new_n_n110_ | new_n_n99_ | new_n_n111_ | new_n_n105_ | new_n_n109_ | new_n_n98_ | new_n_n108_ | new_n_n104_ | new_n_n114_ | new_n_n103_ | new_n_n115_ | new_n_n102_ | new_n_n112_ | new_n_n86_ | new_n_n113_ | new_n_n89_ | new_n_n90_ | new_n_n87_ | new_n_n88_;
  assign new_nv218_ = new_n_n6_ & new_n_n32_;
  assign new_nv229_ = new_n_n2_ & new_n_n18_;
  assign new_n_n9_ = new_n_n123_ | new_n_n124_ | new_n_n125_ | new_n_n126_ | new_n_n129_ | new_n_n127_ | new_n_n128_ | new_n_n138_ | new_n_n149_ | new_n_n139_ | new_n_n133_ | new_n_n148_ | new_n_n132_ | new_n_n142_ | new_n_n131_ | new_n_n143_ | new_n_n137_ | new_n_n141_ | new_n_n130_ | new_n_n140_ | new_n_n136_ | new_n_n146_ | new_n_n135_ | new_n_n147_ | new_n_n134_ | new_n_n144_ | new_n_n118_ | new_n_n145_ | new_n_n121_ | new_n_n122_ | new_n_n119_ | new_n_n120_;
  assign new_nv219_ = new_nv218_ & new_n_n33_;
  assign new_nv228_ = new_nv227_ & new_n_n19_;
  assign new_nv209_ = new_n_n83_ & new_n_n11_ & new_nv207_;
  assign new_n_n5_ = new_n_n41_ | new_n_n42_ | new_n_n39_ | new_n_n40_ | new_n_n45_ | new_n_n43_ | new_n_n49_ | new_n_n44_ | new_n_n47_ | new_n_n48_ | new_n_n34_ | new_n_n46_ | new_n_n37_ | new_n_n38_ | new_n_n35_ | new_n_n36_;
  assign new_nv227_ = new_n_n3_ & new_n_n18_;
  assign new_nv208_ = new_n_n84_ & new_nv207_;
  assign new_nv217_ = new_n_n33_ & new_n_n7_ & new_n_n32_;
  assign new_nv226_ = new_n_n19_ & new_n_n4_ & new_n_n18_;
  assign new_n_n7_ = new_n_n73_ | new_n_n74_ | new_n_n71_ | new_n_n72_ | new_n_n77_ | new_n_n75_ | new_n_n81_ | new_n_n76_ | new_n_n79_ | new_n_n80_ | new_n_n66_ | new_n_n78_ | new_n_n69_ | new_n_n70_ | new_n_n67_ | new_n_n68_;
  assign new_n_n2_ = new_n_n23_ | new_n_n21_ | new_n_n22_ | new_n_n20_;
  assign new_n_n6_ = new_n_n57_ | new_n_n58_ | new_n_n55_ | new_n_n56_ | new_n_n61_ | new_n_n59_ | new_n_n65_ | new_n_n60_ | new_n_n63_ | new_n_n64_ | new_n_n50_ | new_n_n62_ | new_n_n53_ | new_n_n54_ | new_n_n51_ | new_n_n52_;
  assign new_n_n3_ = new_n_n27_ | new_n_n25_ | new_n_n26_ | new_n_n24_;
  assign new_n_n10_ = new_n_n155_ | new_n_n156_ | new_n_n157_ | new_n_n158_ | new_n_n161_ | new_n_n159_ | new_n_n160_ | new_n_n170_ | new_n_n181_ | new_n_n171_ | new_n_n165_ | new_n_n180_ | new_n_n164_ | new_n_n174_ | new_n_n163_ | new_n_n175_ | new_n_n169_ | new_n_n173_ | new_n_n162_ | new_n_n172_ | new_n_n168_ | new_n_n178_ | new_n_n167_ | new_n_n179_ | new_n_n166_ | new_n_n176_ | new_n_n150_ | new_n_n177_ | new_n_n153_ | new_n_n154_ | new_n_n151_ | new_n_n152_;
  assign new_nv212_ = new_n_n83_ & new_n_n9_ & new_n_n85_;
  assign new_n_n4_ = new_n_n31_ | new_n_n29_ | new_n_n30_ | new_n_n28_;
  assign new_n_n11_ = new_n_n187_ | new_n_n188_ | new_n_n189_ | new_n_n190_ | new_n_n193_ | new_n_n191_ | new_n_n192_ | new_n_n202_ | new_n_n213_ | new_n_n203_ | new_n_n197_ | new_n_n212_ | new_n_n196_ | new_n_n206_ | new_n_n195_ | new_n_n207_ | new_n_n201_ | new_n_n205_ | new_n_n194_ | new_n_n204_ | new_n_n200_ | new_n_n210_ | new_n_n199_ | new_n_n211_ | new_n_n198_ | new_n_n208_ | new_n_n182_ | new_n_n209_ | new_n_n185_ | new_n_n186_ | new_n_n183_ | new_n_n184_;
  assign new_nv213_ = new_n_n83_ & new_n_n8_ & new_n_n85_;
  assign new_nv222_ = new_n_n5_ & new_n_n33_;
  assign new_nv210_ = new_n_n83_ & new_n_n10_ & new_nv207_;
  assign new_nv221_ = new_nv220_ & new_n_n33_;
  assign new_nv211_ = new_n_n82_ & new_n_n85_;
  assign new_nv220_ = new_n_n5_ & new_n_n32_;
endmodule


