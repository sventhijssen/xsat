// Benchmark "top" written by ABC on Fri Mar 31 12:12:33 2023

module top ( 
    i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_,
    i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, i_11_,
    i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, i_15_,
    i_32_, i_31_, i_34_, i_33_, i_19_, i_41_, i_36_, i_42_, i_35_, i_43_,
    i_38_, i_29_, i_44_, i_37_,
    o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_,
    o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_,
    o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_,
    o_17_, o_43_, o_30_, o_44_, o_41_, o_42_, o_20_, o_10_, o_9_, o_7_,
    o_8_, o_5_, o_6_, o_3_, o_4_  );
  input  i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_,
    i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_,
    i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_,
    i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_41_, i_36_, i_42_, i_35_,
    i_43_, i_38_, i_29_, i_44_, i_37_;
  output o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_,
    o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_,
    o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_,
    o_17_, o_43_, o_30_, o_44_, o_41_, o_42_, o_20_, o_10_, o_9_, o_7_,
    o_8_, o_5_, o_6_, o_3_, o_4_;
  wire new_ni_40__, new_ni_30__, new_ni_20__, new_ni_9__, new_ni_10__,
    new_ni_7__, new_ni_8__, new_ni_5__, new_ni_6__, new_ni_27__,
    new_ni_14__, new_ni_3__, new_ni_39__, new_ni_28__, new_ni_13__,
    new_ni_4__, new_ni_25__, new_ni_12__, new_ni_1__, new_ni_26__,
    new_ni_11__, new_ni_2__, new_ni_23__, new_ni_18__, new_ni_24__,
    new_ni_17__, new_ni_0__, new_ni_21__, new_ni_16__, new_ni_22__,
    new_ni_15__, new_ni_32__, new_ni_31__, new_ni_34__, new_ni_33__,
    new_ni_19__, new_ni_41__, new_ni_36__, new_ni_42__, new_ni_35__,
    new_ni_43__, new_ni_38__, new_ni_29__, new_ni_44__, new_ni_37__,
    new_no_7__, new_n_n747_, new_n_n736_, new_n_n725_, new_n_n714_,
    new_n_n704_, new_n_n662_, new_n_n651_, new_n_n640_, new_n_n629_,
    new_n_n619_, new_n_n608_, new_n_n598_, new_n_n566_, new_n_n558_,
    new_n_n550_, new_n_n539_, new_n_n530_, new_n_n520_, new_n_n510_,
    new_n_n499_, new_n_n477_, new_n_n467_, new_n_n456_, new_n_n446_,
    new_n_n435_, new_n_n425_, new_n_n414_, new_n_n404_, new_n_n393_,
    new_n_n383_, new_n_n372_, new_n_n362_, new_n_n352_, new_n_n341_,
    new_n_n331_, new_n_n320_, new_n_n310_, new_n_n300_, new_n_n290_,
    new_n_n280_, new_n_n271_, new_n_n264_, new_n_n763_, new_n_n768_,
    new_n_n773_, new_n_n240_, new_n_n235_, new_n_n230_, new_n_n220_,
    new_n_n804_, new_n_n210_, new_n_n205_, new_n_n200_, new_n_n829_,
    new_n_n190_, new_n_n839_, new_n_n856_, new_n_n160_, new_n_n154_,
    new_n_n148_, new_n_n142_, new_n_n879_, new_n_n885_, new_n_n903_,
    new_n_n907_, new_n_n910_, new_n_n84_, new_n_n78_, new_no_41__,
    new_no_23__, new_n_n748_, new_n_n735_, new_n_n726_, new_n_n713_,
    new_n_n705_, new_n_n661_, new_n_n652_, new_n_n639_, new_n_n630_,
    new_n_n618_, new_n_n609_, new_n_n588_, new_n_n565_, new_no_31__,
    new_n_n549_, new_n_n540_, new_no_26__, new_n_n521_, new_n_n509_,
    new_n_n500_, new_n_n476_, new_n_n468_, new_n_n455_, new_n_n447_,
    new_no_18__, new_n_n426_, new_n_n413_, new_n_n405_, new_n_n384_,
    new_n_n382_, new_n_n373_, new_n_n361_, new_no_14__, new_n_n340_,
    new_n_n332_, new_n_n319_, new_n_n311_, new_n_n299_, new_no_10__,
    new_n_n289_, new_no_0__, new_n_n265_, new_n_n258_, new_n_n253_,
    new_n_n246_, new_n_n241_, new_n_n234_, new_n_n788_, new_n_n800_,
    new_n_n803_, new_n_n209_, new_n_n817_, new_n_n199_, new_n_n828_,
    new_n_n835_, new_n_n184_, new_n_n850_, new_n_n860_, new_n_n864_,
    new_n_n870_, new_n_n874_, new_n_n135_, new_n_n131_, new_n_n104_,
    new_n_n98_, new_n_n90_, new_n_n914_, new_n_n77_, new_n_n72_,
    new_no_3__, new_n_n749_, new_n_n734_, new_n_n723_, new_n_n716_,
    new_n_n706_, new_n_n664_, new_n_n653_, new_n_n638_, new_n_n627_,
    new_n_n621_, new_n_n610_, new_n_n579_, new_n_n568_, new_n_n559_,
    new_n_n548_, new_n_n537_, new_n_n531_, new_n_n522_, new_n_n490_,
    new_n_n479_, new_no_22__, new_n_n454_, new_n_n444_, new_n_n437_,
    new_n_n427_, new_n_n412_, new_n_n395_, new_n_n385_, new_n_n360_,
    new_n_n350_, new_n_n343_, new_no_13__, new_n_n318_, new_n_n308_,
    new_n_n302_, new_n_n291_, new_n_n270_, new_n_n263_, new_n_n259_,
    new_n_n254_, new_n_n245_, new_n_n779_, new_n_n782_, new_n_n787_,
    new_n_n801_, new_n_n806_, new_n_n211_, new_n_n816_, new_n_n198_,
    new_n_n830_, new_n_n191_, new_n_n185_, new_n_n851_, new_n_n166_,
    new_n_n155_, new_n_n147_, new_n_n875_, new_n_n878_, new_n_n132_,
    new_n_n118_, new_n_n900_, new_n_n911_, new_n_n915_, new_n_n79_,
    new_n_n923_, new_no_4__, new_n_n750_, new_n_n733_, new_n_n724_,
    new_n_n715_, new_n_n707_, new_n_n663_, new_n_n654_, new_n_n637_,
    new_n_n628_, new_n_n620_, new_n_n611_, new_n_n569_, new_n_n567_,
    new_no_33__, new_n_n547_, new_n_n538_, new_no_27__, new_n_n523_,
    new_n_n489_, new_n_n480_, new_n_n478_, new_no_19__, new_n_n445_,
    new_n_n436_, new_n_n428_, new_n_n403_, new_n_n394_, new_n_n386_,
    new_n_n359_, new_n_n351_, new_n_n342_, new_n_n333_, new_n_n317_,
    new_n_n309_, new_n_n301_, new_n_n292_, new_n_n269_, new_n_n758_,
    new_n_n762_, new_n_n767_, new_n_n774_, new_n_n778_, new_n_n236_,
    new_n_n231_, new_n_n219_, new_n_n805_, new_n_n811_, new_n_n815_,
    new_n_n823_, new_n_n195_, new_n_n834_, new_n_n838_, new_n_n852_,
    new_n_n167_, new_n_n161_, new_n_n871_, new_n_n141_, new_n_n136_,
    new_n_n884_, new_n_n897_, new_n_n111_, new_n_n89_, new_n_n83_,
    new_n_n919_, new_n_n73_, new_n_n754_, new_n_n743_, new_n_n740_,
    new_n_n729_, new_n_n718_, new_n_n708_, new_n_n658_, new_n_n647_,
    new_n_n644_, new_n_n633_, new_n_n623_, new_n_n612_, new_n_n562_,
    new_no_9__, new_n_n553_, new_n_n543_, new_n_n533_, new_n_n524_,
    new_n_n473_, new_n_n463_, new_n_n450_, new_n_n439_, new_n_n429_,
    new_n_n379_, new_n_n368_, new_n_n345_, new_n_n334_, new_n_n286_,
    new_n_n276_, new_n_n255_, new_n_n244_, new_n_n228_, new_n_n796_,
    new_n_n197_, new_n_n831_, new_n_n841_, new_n_n846_, new_n_n146_,
    new_n_n876_, new_n_n881_, new_n_n129_, new_n_n893_, new_n_n88_,
    new_n_n82_, new_n_n75_, new_n_n925_, new_n_n7_, new_n_n753_,
    new_n_n744_, new_n_n739_, new_n_n730_, new_n_n717_, new_n_n709_,
    new_n_n657_, new_n_n648_, new_n_n643_, new_n_n634_, new_n_n622_,
    new_n_n613_, new_no_34__, new_n_n556_, new_n_n552_, new_n_n544_,
    new_n_n532_, new_n_n525_, new_n_n472_, new_n_n464_, new_n_n459_,
    new_n_n438_, new_n_n430_, new_n_n378_, new_n_n369_, new_n_n344_,
    new_n_n335_, new_n_n285_, new_n_n277_, new_n_n761_, new_n_n239_,
    new_n_n790_, new_n_n224_, new_n_n824_, new_n_n194_, new_n_n181_,
    new_n_n176_, new_n_n145_, new_n_n140_, new_n_n887_, new_n_n888_,
    new_n_n124_, new_n_n912_, new_n_n916_, new_n_n921_, new_n_n924_,
    new_no_42__, new_n_n745_, new_n_n738_, new_n_n727_, new_n_n720_,
    new_n_n710_, new_n_n660_, new_n_n649_, new_n_n642_, new_n_n631_,
    new_no_37__, new_n_n614_, new_n_n564_, new_no_30__, new_no_29__,
    new_n_n541_, new_n_n535_, new_n_n526_, new_n_n475_, new_n_n465_,
    new_n_n458_, new_n_n448_, new_n_n431_, new_n_n381_, new_n_n370_,
    new_no_15__, new_n_n353_, new_n_n288_, new_n_n278_, new_n_n757_,
    new_n_n783_, new_n_n229_, new_n_n795_, new_n_n189_, new_n_n840_,
    new_n_n845_, new_n_n144_, new_n_n880_, new_n_n886_, new_n_n913_,
    new_n_n917_, new_n_n920_, new_n_n70_, new_no_43__, new_n_n746_,
    new_n_n737_, new_n_n728_, new_n_n719_, new_n_n711_, new_n_n659_,
    new_n_n650_, new_n_n641_, new_n_n632_, new_n_n624_, new_n_n615_,
    new_n_n563_, new_n_n557_, new_n_n551_, new_n_n542_, new_n_n534_,
    new_n_n527_, new_n_n474_, new_n_n466_, new_n_n457_, new_n_n449_,
    new_n_n440_, new_n_n380_, new_n_n371_, new_n_n363_, new_n_n354_,
    new_n_n287_, new_n_n279_, new_n_n272_, new_n_n789_, new_no_21__,
    new_n_n225_, new_n_n836_, new_n_n183_, new_n_n182_, new_n_n139_,
    new_n_n134_, new_n_n130_, new_n_n87_, new_n_n81_, new_n_n76_,
    new_n_n71_, new_n_n702_, new_n_n691_, new_n_n681_, new_n_n670_,
    new_n_n605_, new_n_n595_, new_n_n584_, new_n_n574_, new_n_n517_,
    new_n_n507_, new_n_n496_, new_n_n485_, new_n_n469_, new_n_n411_,
    new_n_n401_, new_n_n390_, new_n_n375_, new_n_n364_, new_n_n307_,
    new_n_n297_, new_n_n283_, new_n_n273_, new_n_n266_, new_n_n784_,
    new_n_n792_, new_n_n222_, new_n_n215_, new_n_n810_, new_n_n179_,
    new_n_n848_, new_n_n855_, new_n_n859_, new_n_n863_, new_n_n889_,
    new_n_n121_, new_n_n114_, new_n_n902_, new_n_n906_, new_n_n92_,
    new_n_n3_, new_n_n701_, new_n_n692_, new_n_n680_, new_n_n671_,
    new_no_36__, new_n_n596_, new_n_n583_, new_n_n575_, new_no_25__,
    new_n_n508_, new_n_n495_, new_n_n486_, new_n_n460_, new_n_n421_,
    new_n_n400_, new_n_n391_, new_n_n374_, new_n_n365_, new_n_n306_,
    new_n_n298_, new_n_n282_, new_no_6__, new_n_n260_, new_n_n780_,
    new_n_n226_, new_n_n798_, new_n_n214_, new_n_n809_, new_n_n178_,
    new_n_n174_, new_n_n169_, new_n_n163_, new_n_n151_, new_n_n126_,
    new_n_n894_, new_n_n899_, new_n_n107_, new_n_n99_, new_n_n93_,
    new_n_n4_, new_n_n700_, new_no_38__, new_n_n683_, new_n_n672_,
    new_n_n656_, new_n_n604_, new_n_n593_, new_n_n586_, new_n_n576_,
    new_n_n561_, new_n_n554_, new_n_n516_, new_n_n505_, new_n_n498_,
    new_n_n487_, new_n_n471_, new_n_n461_, new_n_n420_, new_n_n410_,
    new_n_n392_, new_n_n377_, new_n_n366_, new_n_n326_, new_n_n316_,
    new_n_n284_, new_n_n274_, new_n_n766_, new_n_n775_, new_n_n791_,
    new_n_n223_, new_n_n814_, new_n_n820_, new_n_n180_, new_n_n847_,
    new_n_n168_, new_n_n157_, new_n_n868_, new_n_n128_, new_n_n122_,
    new_n_n113_, new_n_n105_, new_n_n101_, new_n_n909_, new_n_n5_,
    new_n_n699_, new_n_n690_, new_n_n682_, new_n_n673_, new_n_n646_,
    new_n_n603_, new_n_n594_, new_n_n585_, new_n_n577_, new_n_n560_,
    new_n_n555_, new_n_n515_, new_n_n506_, new_n_n497_, new_n_n488_,
    new_n_n470_, new_n_n462_, new_n_n419_, new_no_17__, new_n_n402_,
    new_n_n376_, new_n_n367_, new_n_n325_, new_no_12__, new_no_8__,
    new_n_n275_, new_n_n771_, new_n_n250_, new_n_n227_, new_n_n797_,
    new_n_n206_, new_n_n202_, new_n_n842_, new_n_n175_, new_n_n162_,
    new_n_n156_, new_n_n867_, new_n_n127_, new_n_n123_, new_n_n112_,
    new_n_n106_, new_n_n100_, new_n_n94_, new_n_n6_, new_n_n698_,
    new_n_n688_, new_n_n677_, new_n_n666_, new_n_n636_, new_n_n602_,
    new_n_n591_, new_n_n580_, new_n_n570_, new_n_n546_, new_no_28__,
    new_n_n514_, new_n_n503_, new_n_n492_, new_n_n481_, new_n_n453_,
    new_n_n442_, new_n_n432_, new_n_n418_, new_n_n408_, new_n_n397_,
    new_no_16__, new_n_n358_, new_n_n348_, new_n_n337_, new_n_n327_,
    new_n_n324_, new_n_n314_, new_n_n304_, new_n_n293_, new_n_n755_,
    new_n_n262_, new_n_n765_, new_n_n251_, new_n_n249_, new_n_n243_,
    new_n_n781_, new_n_n786_, new_n_n218_, new_n_n807_, new_n_n813_,
    new_n_n819_, new_n_n821_, new_n_n826_, new_n_n833_, new_n_n186_,
    new_n_n177_, new_n_n853_, new_n_n165_, new_n_n158_, new_n_n152_,
    new_n_n872_, new_n_n877_, new_n_n133_, new_n_n125_, new_n_n119_,
    new_n_n117_, new_n_n109_, new_n_n904_, new_n_n95_, new_n_n80_,
    new_n_n922_, new_n_n0_, new_n_n697_, new_n_n689_, new_n_n676_,
    new_n_n667_, new_n_n626_, new_n_n601_, new_n_n592_, new_no_35__,
    new_n_n571_, new_n_n545_, new_n_n536_, new_n_n513_, new_n_n504_,
    new_n_n491_, new_n_n482_, new_n_n452_, new_n_n443_, new_n_n422_,
    new_n_n417_, new_n_n409_, new_n_n396_, new_n_n387_, new_n_n357_,
    new_n_n349_, new_n_n336_, new_n_n328_, new_n_n323_, new_n_n315_,
    new_n_n303_, new_n_n294_, new_n_n268_, new_n_n759_, new_n_n256_,
    new_n_n770_, new_n_n772_, new_n_n776_, new_n_n237_, new_n_n232_,
    new_n_n217_, new_n_n213_, new_n_n207_, new_n_n203_, new_no_20__,
    new_n_n825_, new_n_n192_, new_n_n187_, new_n_n172_, new_n_n171_,
    new_n_n857_, new_n_n862_, new_n_n866_, new_n_n150_, new_n_n137_,
    new_n_n883_, new_n_n892_, new_n_n896_, new_n_n116_, new_n_n110_,
    new_n_n905_, new_n_n96_, new_n_n918_, new_n_n74_, new_n_n1_,
    new_n_n696_, new_n_n686_, new_n_n679_, new_n_n668_, new_n_n617_,
    new_n_n600_, new_n_n589_, new_n_n582_, new_n_n572_, new_n_n529_,
    new_n_n518_, new_n_n512_, new_n_n501_, new_n_n494_, new_n_n483_,
    new_n_n451_, new_n_n434_, new_n_n423_, new_n_n416_, new_n_n406_,
    new_n_n399_, new_n_n388_, new_n_n356_, new_n_n346_, new_n_n339_,
    new_n_n329_, new_n_n322_, new_n_n312_, new_no_11__, new_n_n295_,
    new_n_n281_, new_n_n267_, new_n_n261_, new_n_n257_, new_n_n252_,
    new_n_n248_, new_n_n242_, new_no_44__, new_n_n785_, new_n_n793_,
    new_n_n221_, new_n_n802_, new_n_n212_, new_n_n812_, new_n_n204_,
    new_n_n201_, new_n_n196_, new_n_n832_, new_n_n837_, new_n_n843_,
    new_n_n849_, new_n_n854_, new_n_n164_, new_n_n159_, new_n_n153_,
    new_n_n869_, new_n_n143_, new_n_n882_, new_n_n890_, new_n_n120_,
    new_n_n898_, new_n_n901_, new_n_n103_, new_n_n908_, new_no_32__,
    new_n_n85_, new_n_n2_, new_n_n695_, new_n_n687_, new_n_n678_,
    new_n_n669_, new_n_n607_, new_n_n599_, new_n_n590_, new_n_n581_,
    new_n_n573_, new_n_n528_, new_n_n519_, new_n_n511_, new_n_n502_,
    new_n_n493_, new_n_n484_, new_n_n441_, new_n_n433_, new_n_n424_,
    new_n_n415_, new_n_n407_, new_n_n398_, new_n_n389_, new_n_n355_,
    new_n_n347_, new_n_n338_, new_n_n330_, new_n_n321_, new_n_n313_,
    new_n_n305_, new_n_n296_, new_no_5__, new_n_n756_, new_n_n760_,
    new_n_n764_, new_n_n769_, new_n_n247_, new_n_n777_, new_n_n238_,
    new_n_n233_, new_n_n794_, new_n_n799_, new_n_n216_, new_n_n808_,
    new_n_n208_, new_n_n818_, new_n_n822_, new_n_n827_, new_n_n193_,
    new_n_n188_, new_n_n844_, new_n_n173_, new_n_n170_, new_n_n858_,
    new_n_n861_, new_n_n865_, new_n_n149_, new_n_n873_, new_n_n138_,
    new_n_n891_, new_n_n895_, new_n_n115_, new_n_n108_, new_n_n102_,
    new_n_n97_, new_n_n91_, new_n_n86_, new_n_n954_, new_n_n928_,
    new_n_n59_, new_n_n935_, new_n_n938_, new_n_n36_, new_n_n67_,
    new_n_n932_, new_n_n52_, new_n_n43_, new_n_n37_, new_n_n68_,
    new_n_n58_, new_n_n50_, new_n_n45_, new_n_n38_, new_n_n927_,
    new_n_n57_, new_n_n51_, new_n_n44_, new_n_n941_, new_n_n955_,
    new_n_n685_, new_n_n674_, new_n_n578_, new_n_n69_, new_n_n32_,
    new_n_n947_, new_n_n15_, new_n_n8_, new_n_n684_, new_n_n675_,
    new_n_n587_, new_n_n926_, new_n_n31_, new_n_n24_, new_n_n950_,
    new_n_n953_, new_n_n703_, new_n_n693_, new_n_n597_, new_n_n945_,
    new_n_n22_, new_n_n17_, new_n_n9_, new_no_39__, new_n_n694_,
    new_n_n606_, new_n_n30_, new_n_n23_, new_n_n16_, new_n_n10_,
    new_n_n722_, new_no_40__, new_n_n616_, new_n_n49_, new_n_n939_,
    new_n_n943_, new_n_n27_, new_n_n18_, new_n_n952_, new_n_n721_,
    new_n_n712_, new_n_n625_, new_n_n936_, new_n_n42_, new_n_n34_,
    new_n_n946_, new_n_n949_, new_n_n11_, new_n_n742_, new_n_n731_,
    new_n_n635_, new_n_n63_, new_n_n933_, new_n_n33_, new_n_n25_,
    new_n_n20_, new_n_n12_, new_n_n741_, new_n_n732_, new_n_n645_,
    new_n_n62_, new_n_n56_, new_n_n944_, new_n_n26_, new_n_n19_,
    new_n_n13_, new_n_n751_, new_n_n655_, new_n_n929_, new_n_n930_,
    new_n_n54_, new_n_n46_, new_n_n39_, new_n_n948_, new_n_n951_,
    new_no_1__, new_n_n752_, new_n_n665_, new_n_n64_, new_n_n61_,
    new_n_n55_, new_n_n937_, new_n_n940_, new_n_n21_, new_n_n14_,
    new_n_n65_, new_n_n60_, new_n_n53_, new_n_n48_, new_n_n40_,
    new_n_n942_, new_n_n28_, new_n_n66_, new_n_n931_, new_n_n934_,
    new_n_n47_, new_n_n41_, new_n_n35_, new_n_n29_;
  assign o_1_ = new_no_1__;
  assign o_19_ = new_no_19__;
  assign o_2_ = new_no_42__;
  assign o_0_ = new_no_0__;
  assign new_ni_40__ = i_40_;
  assign o_29_ = new_no_29__;
  assign new_ni_30__ = i_30_;
  assign o_39_ = new_no_39__;
  assign o_38_ = new_no_38__;
  assign o_25_ = new_no_25__;
  assign o_12_ = new_no_12__;
  assign o_37_ = new_no_37__;
  assign o_26_ = new_no_26__;
  assign o_11_ = new_no_11__;
  assign new_ni_20__ = i_20_;
  assign o_36_ = new_no_36__;
  assign o_27_ = new_no_27__;
  assign o_14_ = new_no_14__;
  assign new_ni_9__ = i_9_;
  assign o_35_ = new_no_35__;
  assign o_28_ = new_no_28__;
  assign o_13_ = new_no_13__;
  assign o_34_ = new_no_34__;
  assign o_21_ = new_no_21__;
  assign o_16_ = new_no_16__;
  assign new_ni_10__ = i_10_;
  assign new_ni_7__ = i_7_;
  assign o_40_ = new_no_40__;
  assign o_33_ = new_no_33__;
  assign o_22_ = new_no_22__;
  assign o_15_ = new_no_15__;
  assign new_ni_8__ = i_8_;
  assign o_32_ = new_no_32__;
  assign o_23_ = new_no_23__;
  assign o_18_ = new_no_18__;
  assign new_ni_5__ = i_5_;
  assign o_31_ = new_no_31__;
  assign o_24_ = new_no_44__;
  assign o_17_ = new_no_17__;
  assign new_ni_6__ = i_6_;
  assign o_43_ = new_no_43__;
  assign o_30_ = new_no_30__;
  assign new_ni_27__ = i_27_;
  assign new_ni_14__ = i_14_;
  assign new_ni_3__ = i_3_;
  assign o_44_ = new_no_44__;
  assign new_ni_39__ = i_39_;
  assign new_ni_28__ = i_28_;
  assign new_ni_13__ = i_13_;
  assign new_ni_4__ = i_4_;
  assign o_41_ = new_no_41__;
  assign new_ni_25__ = i_25_;
  assign new_ni_12__ = i_12_;
  assign new_ni_1__ = i_1_;
  assign o_42_ = new_no_42__;
  assign o_20_ = new_no_20__;
  assign new_ni_26__ = i_26_;
  assign new_ni_11__ = i_11_;
  assign new_ni_2__ = i_2_;
  assign new_ni_23__ = i_23_;
  assign new_ni_18__ = i_18_;
  assign new_ni_24__ = i_24_;
  assign new_ni_17__ = i_17_;
  assign new_ni_0__ = i_0_;
  assign o_10_ = new_no_10__;
  assign new_ni_21__ = i_21_;
  assign new_ni_16__ = i_16_;
  assign new_ni_22__ = i_22_;
  assign new_ni_15__ = i_15_;
  assign o_9_ = new_no_9__;
  assign new_ni_32__ = i_32_;
  assign new_ni_31__ = i_31_;
  assign o_7_ = new_no_7__;
  assign new_ni_34__ = i_34_;
  assign o_8_ = new_no_8__;
  assign new_ni_33__ = i_33_;
  assign new_ni_19__ = i_19_;
  assign o_5_ = new_no_5__;
  assign new_ni_41__ = i_41_;
  assign new_ni_36__ = i_36_;
  assign o_6_ = new_no_6__;
  assign new_ni_42__ = i_42_;
  assign new_ni_35__ = i_35_;
  assign o_3_ = new_no_3__;
  assign new_ni_43__ = i_43_;
  assign new_ni_38__ = i_38_;
  assign new_ni_29__ = i_29_;
  assign o_4_ = new_no_4__;
  assign new_ni_44__ = i_44_;
  assign new_ni_37__ = i_37_;
  assign new_no_7__ = new_n_n877_ | new_n_n898_ | new_n_n932_;
  assign new_n_n747_ = ~new_ni_29__;
  assign new_n_n736_ = ~new_ni_16__;
  assign new_n_n725_ = ~new_ni_12__;
  assign new_n_n714_ = ~new_ni_44__;
  assign new_n_n704_ = new_n_n709_ | new_n_n708_ | new_n_n707_;
  assign new_n_n662_ = new_n_n869_ | new_n_n871_ | new_n_n872_;
  assign new_n_n651_ = new_n_n930_ | new_n_n931_ | new_n_n932_;
  assign new_n_n640_ = new_n_n672_ | new_n_n671_ | new_n_n670_;
  assign new_n_n629_ = new_n_n640_ | new_n_n639_ | new_n_n638_;
  assign new_n_n619_ = new_n_n853_ | new_n_n854_ | new_n_n860_;
  assign new_n_n608_ = new_n_n617_ | new_n_n616_ | new_n_n615_;
  assign new_n_n598_ = new_n_n804_ | new_n_n808_ | new_n_n819_;
  assign new_n_n566_ = new_n_n577_ | new_n_n576_ | new_n_n575_;
  assign new_n_n558_ = new_n_n853_ | new_n_n867_ | new_n_n898_;
  assign new_n_n550_ = new_no_44__ | new_n_n788_ | new_n_n789_;
  assign new_n_n539_ = new_n_n548_ | new_n_n547_ | new_n_n546_;
  assign new_n_n530_ = new_n_n774_ | new_n_n780_ | new_n_n792_;
  assign new_n_n520_ = new_n_n529_ | new_n_n528_ | new_n_n527_;
  assign new_n_n510_ = new_n_n790_ | new_n_n791_ | new_n_n792_;
  assign new_n_n499_ = new_n_n826_ | new_n_n827_ | new_n_n830_;
  assign new_n_n477_ = new_n_n495_ | new_n_n494_ | new_n_n493_;
  assign new_n_n467_ = new_n_n779_ | new_n_n780_ | new_no_44__;
  assign new_n_n456_ = new_n_n576_ | new_n_n461_ | new_n_n460_;
  assign new_n_n446_ = new_n_n800_ | new_n_n803_ | new_n_n804_;
  assign new_n_n435_ = new_n_n437_ | new_n_n438_;
  assign new_n_n425_ = new_n_n805_ | new_n_n808_ | new_n_n817_;
  assign new_n_n414_ = new_n_n423_ | new_n_n422_ | new_n_n311_;
  assign new_n_n404_ = new_n_n802_ | new_n_n805_ | new_n_n807_;
  assign new_n_n393_ = new_n_n407_ | new_n_n406_ | new_n_n405_;
  assign new_n_n383_ = new_n_n782_ | new_n_n783_ | new_n_n785_;
  assign new_n_n372_ = new_n_n889_ | new_n_n945_ | new_n_n948_;
  assign new_n_n362_ = new_n_n778_ | new_no_21__ | new_n_n791_;
  assign new_n_n352_ = new_n_n767_ | new_n_n768_ | new_n_n770_;
  assign new_n_n341_ = new_n_n824_ | new_n_n826_ | new_n_n833_;
  assign new_n_n331_ = new_n_n781_ | new_n_n783_ | new_n_n784_;
  assign new_n_n320_ = new_n_n328_ | new_n_n327_ | new_n_n326_;
  assign new_n_n310_ = new_n_n836_ | new_n_n841_ | new_n_n953_;
  assign new_n_n300_ = new_n_n808_ | new_n_n810_ | new_n_n814_;
  assign new_n_n290_ = new_n_n843_ | new_n_n853_ | new_n_n867_;
  assign new_n_n280_ = new_n_n879_ | new_n_n882_ | new_n_n889_;
  assign new_n_n271_ = new_n_n884_ | new_n_n891_ | new_n_n896_;
  assign new_n_n264_ = new_n_n750_ & new_ni_29__ & new_ni_30__;
  assign new_n_n763_ = new_n_n185_ & new_n_n260_ & new_ni_30__;
  assign new_n_n768_ = new_n_n254_ & new_n_n253_ & new_ni_30__;
  assign new_n_n773_ = new_n_n247_ & new_n_n248_;
  assign new_n_n240_ = new_ni_30__ & new_ni_29__;
  assign new_n_n235_ = new_ni_21__ & new_ni_25__ & new_n_n750_;
  assign new_n_n230_ = new_ni_21__ & new_ni_22__ & new_ni_28__;
  assign new_n_n220_ = new_ni_20__ & new_n_n751_ & new_ni_27__;
  assign new_n_n804_ = new_n_n143_ & new_n_n133_ & new_n_n232_;
  assign new_n_n210_ = new_ni_18__ & new_ni_19__ & new_ni_21__;
  assign new_n_n205_ = new_n_n751_ & new_ni_22__ & new_ni_30__;
  assign new_n_n200_ = new_n_n741_ & new_n_n754_ & new_ni_19__;
  assign new_n_n829_ = new_n_n270_ & new_n_n84_ & new_ni_30__;
  assign new_n_n190_ = new_ni_24__ & new_n_n750_ & new_n_n747_;
  assign new_n_n839_ = new_n_n185_ & new_n_n184_ & new_n_n753_;
  assign new_n_n856_ = new_n_n169_ & new_n_n168_ & new_ni_31__;
  assign new_n_n160_ = new_ni_27__ & new_n_n747_ & new_n_n753_;
  assign new_n_n154_ = new_ni_8__ & new_ni_16__ & new_ni_18__;
  assign new_n_n148_ = new_n_n749_ & new_n_n751_ & new_ni_25__;
  assign new_n_n142_ = new_ni_13__ & new_n_n739_ & new_n_n751_;
  assign new_n_n879_ = new_n_n192_ & new_n_n136_ & new_n_n217_;
  assign new_n_n885_ = new_ni_30__ & new_n_n131_;
  assign new_n_n903_ = new_n_n753_ & new_n_n105_;
  assign new_n_n907_ = new_n_n753_ & new_n_n98_;
  assign new_n_n910_ = new_n_n107_ & new_n_n91_ & new_n_n234_;
  assign new_n_n84_ = new_ni_26__ & new_n_n750_ & new_n_n747_;
  assign new_n_n78_ = new_ni_0__ & new_n_n745_ & new_n_n754_;
  assign new_no_41__ = new_n_n232_ & new_n_n72_;
  assign new_no_23__ = new_n_n764_ | new_n_n759_;
  assign new_n_n748_ = ~new_ni_26__;
  assign new_n_n735_ = ~new_ni_0__;
  assign new_n_n726_ = ~new_ni_4__;
  assign new_n_n713_ = ~new_ni_43__;
  assign new_n_n705_ = new_n_n847_ | new_n_n851_ | new_n_n859_;
  assign new_n_n661_ = new_n_n874_ | new_n_n875_ | new_n_n876_;
  assign new_n_n652_ = new_n_n915_ | new_n_n917_ | new_no_41__;
  assign new_n_n639_ = new_n_n669_ | new_n_n668_ | new_n_n667_;
  assign new_n_n630_ = new_n_n643_ | new_n_n642_ | new_n_n641_;
  assign new_n_n618_ = new_n_n861_ | new_n_n862_ | new_n_n867_;
  assign new_n_n609_ = new_n_n620_ | new_n_n619_ | new_n_n618_;
  assign new_n_n588_ = new_n_n603_ | new_n_n602_ | new_n_n601_;
  assign new_n_n565_ = new_n_n574_ | new_n_n573_ | new_n_n572_;
  assign new_no_31__ = new_n_n909_ | new_n_n559_;
  assign new_n_n549_ = new_n_n793_ | new_n_n796_ | new_n_n799_;
  assign new_n_n540_ = new_n_n551_ | new_n_n550_ | new_n_n549_;
  assign new_no_26__ = new_n_n794_ | new_n_n530_;
  assign new_n_n521_ = new_n_n846_ | new_n_n855_ | new_n_n876_;
  assign new_n_n509_ = new_n_n793_ | new_n_n794_ | new_n_n795_;
  assign new_n_n500_ = new_n_n823_ | new_n_n824_ | new_n_n825_;
  assign new_n_n476_ = new_n_n492_ | new_n_n491_ | new_n_n490_;
  assign new_n_n468_ = new_n_n769_ | new_n_n774_ | new_n_n775_;
  assign new_n_n455_ = new_n_n486_ | new_n_n459_ | new_n_n458_;
  assign new_n_n447_ = new_n_n792_ | new_n_n794_ | new_n_n796_;
  assign new_no_18__ = new_n_n435_ | new_n_n436_;
  assign new_n_n426_ = new_n_n799_ | new_n_n802_ | new_n_n803_;
  assign new_n_n413_ = new_n_n421_ | new_n_n420_ | new_n_n419_;
  assign new_n_n405_ = new_n_n797_ | new_n_n800_ | new_n_n801_;
  assign new_n_n384_ = new_n_n776_ | new_n_n777_ | new_n_n778_;
  assign new_n_n382_ = new_n_n786_ | new_n_n789_ | new_no_21__;
  assign new_n_n373_ = new_n_n872_ | new_n_n885_ | new_n_n886_;
  assign new_n_n361_ = new_n_n795_ | new_n_n798_ | new_n_n799_;
  assign new_no_14__ = new_n_n949_ | new_n_n353_;
  assign new_n_n340_ = new_n_n855_ | new_n_n870_ | new_n_n937_;
  assign new_n_n332_ = new_n_n769_ | new_n_n770_ | new_n_n771_;
  assign new_n_n319_ = new_n_n325_ | new_n_n324_ | new_n_n323_;
  assign new_n_n311_ = new_n_n827_ | new_n_n830_ | new_n_n831_;
  assign new_n_n299_ = new_n_n817_ | new_no_20__ | new_n_n827_;
  assign new_no_10__ = new_n_n291_ | new_n_n292_;
  assign new_n_n289_ = new_n_n889_ | new_n_n903_ | new_n_n906_;
  assign new_no_0__ = new_n_n271_ | new_n_n272_;
  assign new_n_n265_ = new_n_n754_ & new_n_n752_ & new_n_n751_;
  assign new_n_n258_ = new_n_n752_ & new_ni_20__ & new_ni_21__;
  assign new_n_n253_ = new_n_n751_ & new_ni_22__ & new_n_n747_;
  assign new_n_n246_ = new_n_n754_ & new_n_n752_ & new_n_n749_;
  assign new_n_n241_ = new_n_n751_ & new_ni_22__ & new_ni_28__;
  assign new_n_n234_ = new_n_n753_ & new_ni_29__;
  assign new_n_n788_ = new_n_n206_ & new_n_n250_;
  assign new_n_n800_ = new_n_n221_ & new_n_n220_ & new_n_n247_;
  assign new_n_n803_ = new_n_n216_ & new_n_n215_ & new_n_n214_;
  assign new_n_n209_ = new_ni_30__ & new_ni_26__;
  assign new_n_n817_ = new_n_n195_ & new_n_n25_ & new_n_n240_;
  assign new_n_n199_ = new_ni_20__ & new_n_n751_ & new_ni_22__;
  assign new_n_n828_ = new_n_n263_ & new_n_n196_ & new_ni_30__;
  assign new_n_n835_ = new_n_n270_ & new_n_n190_ & new_ni_30__;
  assign new_n_n184_ = new_ni_22__ & new_ni_28__ & new_n_n747_;
  assign new_n_n850_ = new_n_n179_ & new_n_n172_ & new_n_n232_;
  assign new_n_n860_ = new_n_n162_ & new_n_n161_ & new_n_n160_;
  assign new_n_n864_ = new_n_n263_ & new_n_n155_ & new_n_n753_;
  assign new_n_n870_ = new_n_n149_ & new_n_n148_ & new_n_n232_;
  assign new_n_n874_ = new_n_n143_ & new_n_n203_ & new_n_n198_;
  assign new_n_n135_ = new_ni_5__ & new_n_n754_ & new_ni_19__;
  assign new_n_n131_ = new_n_n132_ & new_n_n161_ & new_n_n184_;
  assign new_n_n104_ = new_ni_0__ & new_n_n743_ & new_n_n727_;
  assign new_n_n98_ = new_n_n99_ & new_n_n166_ & new_n_n257_;
  assign new_n_n90_ = new_n_n738_ & new_ni_16__ & new_n_n754_;
  assign new_n_n914_ = new_ni_30__ & new_n_n85_;
  assign new_n_n77_ = new_ni_26__ & new_n_n747_ & new_ni_30__;
  assign new_n_n72_ = new_n_n101_ & new_n_n242_ & new_n_n223_;
  assign new_no_3__ = new_n_n854_ | new_n_n829_;
  assign new_n_n749_ = ~new_ni_20__;
  assign new_n_n734_ = ~new_ni_31__;
  assign new_n_n723_ = ~new_ni_33__;
  assign new_n_n716_ = ~new_ni_36__;
  assign new_n_n706_ = new_n_n810_ | new_n_n814_ | new_no_20__;
  assign new_n_n664_ = new_n_n862_ | new_n_n863_ | new_n_n865_;
  assign new_n_n653_ = new_n_n911_ | new_n_n912_ | new_n_n914_;
  assign new_n_n638_ = new_n_n666_ | new_n_n665_ | new_n_n664_;
  assign new_n_n627_ = new_n_n634_ | new_n_n633_ | new_n_n955_;
  assign new_n_n621_ = new_n_n822_ | new_n_n826_ | new_n_n829_;
  assign new_n_n610_ = new_n_n623_ | new_n_n622_ | new_n_n621_;
  assign new_n_n579_ = new_n_n755_ | new_n_n758_ | new_n_n763_;
  assign new_n_n568_ = new_n_n949_ | new_n_n953_ | new_n_n955_;
  assign new_n_n559_ = new_n_n867_ | new_n_n874_ | new_n_n882_;
  assign new_n_n548_ = new_n_n807_ | new_n_n811_ | new_n_n815_;
  assign new_n_n537_ = new_n_n541_ | new_n_n542_;
  assign new_n_n531_ = new_n_n535_ | new_n_n534_ | new_n_n533_;
  assign new_n_n522_ = new_n_n828_ | new_n_n833_ | new_n_n842_;
  assign new_n_n490_ = new_n_n904_ | new_n_n908_ | new_n_n937_;
  assign new_n_n479_ = new_n_n501_ | new_n_n500_ | new_n_n499_;
  assign new_no_22__ = new_n_n469_ | new_n_n470_;
  assign new_n_n454_ = new_n_n457_ | new_n_n456_ | new_n_n953_;
  assign new_n_n444_ = new_n_n833_ | new_n_n855_ | new_n_n864_;
  assign new_n_n437_ = new_n_n442_ | new_n_n443_;
  assign new_n_n427_ = new_n_n795_ | new_n_n796_ | new_n_n798_;
  assign new_n_n412_ = new_n_n486_ | new_n_n418_ | new_n_n417_;
  assign new_n_n395_ = new_n_n955_ | new_n_n944_;
  assign new_n_n385_ = new_n_n769_ | new_n_n772_ | new_n_n773_;
  assign new_n_n360_ = new_n_n800_ | new_n_n801_ | new_n_n802_;
  assign new_n_n350_ = new_n_n775_ | new_n_n776_ | new_n_n778_;
  assign new_n_n343_ = new_n_n814_ | new_n_n816_ | new_n_n819_;
  assign new_no_13__ = new_n_n333_ | new_n_n334_;
  assign new_n_n318_ = new_n_n486_ | new_n_n322_ | new_n_n321_;
  assign new_n_n308_ = new_n_n314_ | new_n_n313_ | new_n_n312_;
  assign new_n_n302_ = new_n_n795_ | new_n_n797_ | new_n_n801_;
  assign new_n_n291_ = new_n_n293_ | new_n_n294_;
  assign new_n_n270_ = new_n_n754_ & new_ni_19__ & new_ni_21__;
  assign new_n_n263_ = new_n_n754_ & new_n_n752_ & new_ni_20__;
  assign new_n_n259_ = new_ni_21__ & new_n_n748_ & new_ni_29__;
  assign new_n_n254_ = new_n_n754_ & new_ni_19__ & new_n_n749_;
  assign new_n_n245_ = new_n_n751_ & new_n_n750_ & new_n_n747_;
  assign new_n_n779_ = new_n_n250_ & new_n_n253_ & new_ni_30__;
  assign new_n_n782_ = new_n_n246_ & new_n_n237_ & new_ni_30__;
  assign new_n_n787_ = new_n_n254_ & new_n_n231_ & new_ni_30__;
  assign new_n_n801_ = new_n_n246_ & new_n_n223_ & new_n_n240_;
  assign new_n_n806_ = new_n_n262_ & new_n_n224_ & new_n_n753_;
  assign new_n_n211_ = new_n_n743_ & new_n_n754_ & new_n_n752_;
  assign new_n_n816_ = new_n_n242_ & new_n_n233_ & new_n_n232_;
  assign new_n_n198_ = new_ni_28__ & new_n_n747_ & new_ni_30__;
  assign new_n_n830_ = new_n_n195_ & new_n_n235_ & new_n_n240_;
  assign new_n_n191_ = new_ni_20__ & new_ni_21__ & new_n_n747_;
  assign new_n_n185_ = new_n_n754_ & new_ni_20__ & new_n_n751_;
  assign new_n_n851_ = new_n_n135_ & new_n_n199_ & new_n_n217_;
  assign new_n_n166_ = new_n_n752_ & new_ni_20__ & new_n_n751_;
  assign new_n_n155_ = new_ni_21__ & new_ni_24__ & new_ni_29__;
  assign new_n_n147_ = new_n_n750_ & new_ni_29__ & new_ni_38__;
  assign new_n_n875_ = new_n_n142_ & new_n_n141_ & new_n_n753_;
  assign new_n_n878_ = new_n_n137_ & new_n_n148_ & new_ni_30__;
  assign new_n_n132_ = new_ni_2__ & new_n_n744_ & new_n_n754_;
  assign new_n_n118_ = new_n_n183_ & new_n_n215_ & new_n_n119_;
  assign new_n_n900_ = new_n_n113_ & new_n_n112_ & new_n_n111_;
  assign new_n_n911_ = new_n_n90_ & new_n_n88_ & new_n_n208_;
  assign new_n_n915_ = new_ni_30__ & new_n_n83_;
  assign new_n_n79_ = new_n_n735_ & new_ni_18__ & new_n_n752_;
  assign new_n_n923_ = new_n_n73_ & new_n_n199_ & new_n_n269_;
  assign new_no_4__ = new_n_n829_ | new_n_n835_ | new_n_n896_;
  assign new_n_n750_ = ~new_ni_28__;
  assign new_n_n733_ = ~new_ni_5__;
  assign new_n_n724_ = ~new_ni_13__;
  assign new_n_n715_ = ~new_ni_40__;
  assign new_n_n707_ = new_n_n803_ | new_n_n805_ | new_n_n808_;
  assign new_n_n663_ = new_n_n866_ | new_n_n867_ | new_n_n868_;
  assign new_n_n654_ = new_n_n907_ | new_n_n909_ | new_no_32__;
  assign new_n_n637_ = new_n_n663_ | new_n_n662_ | new_n_n661_;
  assign new_n_n628_ = new_n_n637_ | new_n_n636_ | new_n_n635_;
  assign new_n_n620_ = new_n_n835_ | new_n_n839_ | new_n_n841_;
  assign new_n_n611_ = new_n_n711_ | new_n_n710_ | new_n_n624_;
  assign new_n_n569_ = new_n_n917_ | new_n_n941_ | new_n_n943_;
  assign new_n_n567_ = new_n_n579_ | new_n_n578_ | new_n_n314_;
  assign new_no_33__ = new_n_n560_ | new_n_n561_;
  assign new_n_n547_ = new_n_n817_ | new_n_n818_ | new_n_n821_;
  assign new_n_n538_ = new_n_n545_ | new_n_n544_ | new_n_n543_;
  assign new_no_27__ = new_n_n532_ | new_n_n531_;
  assign new_n_n523_ = new_n_n816_ | new_n_n818_ | new_n_n819_;
  assign new_n_n489_ = new_n_n945_ | new_n_n948_ | new_n_n949_;
  assign new_n_n480_ = new_n_n504_ | new_n_n503_ | new_n_n502_;
  assign new_n_n478_ = new_n_n498_ | new_n_n497_ | new_n_n496_;
  assign new_no_19__ = new_n_n454_ | new_n_n455_;
  assign new_n_n445_ = new_n_n816_ | new_n_n820_ | new_n_n827_;
  assign new_n_n436_ = new_n_n441_ | new_n_n440_ | new_n_n439_;
  assign new_n_n428_ = new_no_21__ | new_n_n790_ | new_n_n791_;
  assign new_n_n403_ = new_n_n810_ | new_n_n814_ | new_n_n816_;
  assign new_n_n394_ = new_n_n410_ | new_n_n409_ | new_n_n408_;
  assign new_n_n386_ = new_n_n764_ | new_n_n766_ | new_n_n768_;
  assign new_n_n359_ = new_n_n814_ | new_n_n817_ | new_no_20__;
  assign new_n_n351_ = new_n_n772_ | new_n_n773_ | new_n_n774_;
  assign new_n_n342_ = new_n_n821_ | new_no_20__ | new_n_n823_;
  assign new_n_n333_ = new_n_n335_ | new_n_n336_;
  assign new_n_n317_ = new_n_n320_ | new_n_n319_ | new_n_n955_;
  assign new_n_n309_ = new_n_n687_ | new_n_n316_ | new_n_n315_;
  assign new_n_n301_ = new_n_n802_ | new_n_n803_ | new_n_n805_;
  assign new_n_n292_ = new_n_n486_ | new_n_n296_ | new_n_n295_;
  assign new_n_n269_ = new_ni_28__ & new_ni_29__ & new_n_n753_;
  assign new_n_n758_ = new_n_n264_ & new_n_n265_;
  assign new_n_n762_ = new_n_n263_ & new_n_n259_ & new_n_n753_;
  assign new_n_n767_ = new_n_n205_ & new_n_n255_;
  assign new_n_n774_ = new_n_n246_ & new_n_n245_ & new_ni_30__;
  assign new_n_n778_ = new_n_n242_ & new_n_n241_ & new_n_n240_;
  assign new_n_n236_ = new_n_n745_ & new_ni_18__ & new_ni_20__;
  assign new_n_n231_ = new_n_n751_ & new_ni_23__ & new_n_n747_;
  assign new_n_n219_ = new_ni_11__ & new_ni_18__ & new_n_n752_;
  assign new_n_n805_ = new_n_n250_ & new_n_n229_ & new_n_n234_;
  assign new_n_n811_ = new_n_n218_ & new_n_n211_;
  assign new_n_n815_ = new_n_n206_ & new_n_n268_;
  assign new_n_n823_ = new_n_n200_ & new_n_n199_ & new_n_n198_;
  assign new_n_n195_ = new_ni_11__ & new_n_n752_ & new_ni_20__;
  assign new_n_n834_ = new_n_n192_ & new_n_n191_ & new_ni_30__;
  assign new_n_n838_ = new_n_n187_ & new_n_n186_ & new_n_n234_;
  assign new_n_n852_ = new_n_n268_ & new_n_n225_ & new_n_n232_;
  assign new_n_n167_ = new_n_n741_ & new_ni_6__ & new_n_n754_;
  assign new_n_n161_ = new_ni_19__ & new_ni_20__ & new_n_n751_;
  assign new_n_n871_ = new_n_n183_ & new_n_n215_ & new_n_n147_;
  assign new_n_n141_ = new_n_n746_ & new_n_n750_ & new_n_n747_;
  assign new_n_n136_ = new_n_n749_ & new_n_n751_ & new_ni_26__;
  assign new_n_n884_ = new_n_n79_ & new_n_n133_ & new_n_n232_;
  assign new_n_n897_ = new_ni_41__ & new_n_n118_;
  assign new_n_n111_ = new_n_n750_ & new_n_n747_ & new_n_n753_;
  assign new_n_n89_ = new_n_n737_ & new_n_n736_ & new_n_n754_;
  assign new_n_n83_ = new_n_n101_ & new_n_n258_ & new_n_n84_;
  assign new_n_n919_ = new_n_n79_ & new_n_n203_ & new_n_n217_;
  assign new_n_n73_ = new_n_n735_ & new_n_n754_ & new_ni_19__;
  assign new_n_n754_ = ~new_ni_18__;
  assign new_n_n743_ = ~new_ni_10__;
  assign new_n_n740_ = ~new_ni_9__;
  assign new_n_n729_ = ~new_ni_23__;
  assign new_n_n718_ = ~new_ni_34__;
  assign new_n_n708_ = new_n_n783_ | new_no_21__ | new_n_n802_;
  assign new_n_n658_ = new_n_n890_ | new_n_n892_ | new_n_n893_;
  assign new_n_n647_ = new_n_n685_ | new_n_n384_ | new_n_n467_;
  assign new_n_n644_ = new_n_n680_ | new_n_n506_ | new_n_n505_;
  assign new_n_n633_ = new_n_n651_ | new_n_n650_ | new_n_n649_;
  assign new_n_n623_ = new_n_n791_ | new_n_n797_ | new_n_n800_;
  assign new_n_n612_ = new_n_n914_ | new_n_n928_ | new_n_n944_;
  assign new_n_n562_ = new_n_n568_ | new_n_n564_;
  assign new_no_9__ = new_n_n860_ | new_n_n868_ | new_n_n872_;
  assign new_n_n553_ = new_n_n273_ | new_n_n556_ | new_no_9__;
  assign new_n_n543_ = new_n_n876_ | new_n_n880_ | new_n_n890_;
  assign new_n_n533_ = new_n_n859_ | new_n_n860_ | new_n_n872_;
  assign new_n_n524_ = new_n_n809_ | new_n_n811_ | new_n_n815_;
  assign new_n_n473_ = new_n_n483_ | new_n_n482_ | new_n_n481_;
  assign new_n_n463_ = new_n_n804_ | new_n_n807_ | new_n_n808_;
  assign new_n_n450_ = new_n_n773_ | new_n_n774_ | new_n_n777_;
  assign new_n_n439_ = new_n_n448_ | new_n_n447_ | new_n_n446_;
  assign new_n_n429_ = new_n_n786_ | new_n_n788_ | new_n_n789_;
  assign new_n_n379_ = new_n_n806_ | new_n_n808_ | new_n_n810_;
  assign new_n_n368_ = new_n_n380_ | new_n_n379_ | new_n_n378_;
  assign new_n_n345_ = new_n_n801_ | new_n_n802_ | new_n_n803_;
  assign new_n_n334_ = new_n_n339_ | new_n_n338_ | new_n_n337_;
  assign new_n_n286_ = new_n_n946_ | new_n_n947_ | new_n_n950_;
  assign new_n_n276_ = new_n_n283_ | new_n_n282_ | new_n_n281_;
  assign new_n_n255_ = new_ni_18__ & new_n_n752_ & new_ni_20__;
  assign new_n_n244_ = new_n_n751_ & new_ni_23__ & new_ni_30__;
  assign new_n_n228_ = new_n_n751_ & new_ni_23__ & new_n_n750_;
  assign new_n_n796_ = new_n_n262_ & new_n_n224_ & new_ni_30__;
  assign new_n_n197_ = new_ni_3__ & new_n_n754_ & new_ni_19__;
  assign new_n_n831_ = new_n_n254_ & new_n_n194_ & new_n_n234_;
  assign new_n_n841_ = new_n_n182_ & new_n_n218_ & new_n_n264_;
  assign new_n_n846_ = new_n_n176_ & new_n_n235_ & new_n_n232_;
  assign new_n_n146_ = new_ni_0__ & new_ni_2__ & new_n_n744_;
  assign new_n_n876_ = new_n_n140_ & new_n_n218_ & new_n_n214_;
  assign new_n_n881_ = new_n_n134_ & new_n_n178_ & new_n_n232_;
  assign new_n_n129_ = new_n_n733_ & new_ni_15__ & new_ni_18__;
  assign new_n_n893_ = new_n_n124_ & new_n_n166_ & new_n_n198_;
  assign new_n_n88_ = new_ni_19__ & new_ni_20__ & new_ni_22__;
  assign new_n_n82_ = new_ni_0__ & new_n_n733_ & new_ni_18__;
  assign new_n_n75_ = new_n_n747_ & new_ni_27__;
  assign new_n_n925_ = new_n_n120_ & new_n_n136_ & new_n_n198_;
  assign new_n_n7_ = new_ni_29__ & new_n_n753_ & new_n_n730_;
  assign new_n_n753_ = ~new_ni_30__;
  assign new_n_n744_ = ~new_ni_3__;
  assign new_n_n739_ = ~new_ni_14__;
  assign new_n_n730_ = ~new_ni_38__;
  assign new_n_n717_ = ~new_ni_35__;
  assign new_n_n709_ = new_n_n769_ | new_n_n772_ | new_n_n776_;
  assign new_n_n657_ = new_n_n894_ | new_n_n897_ | new_n_n898_;
  assign new_n_n648_ = new_n_n687_ | new_n_n451_ | new_n_n686_;
  assign new_n_n643_ = new_n_n504_ | new_n_n679_ | new_n_n678_;
  assign new_n_n634_ = new_n_n654_ | new_n_n653_ | new_n_n652_;
  assign new_n_n622_ = new_n_n802_ | new_n_n806_ | new_n_n813_;
  assign new_n_n613_ = new_no_32__ | new_n_n911_ | new_n_n912_;
  assign new_no_34__ = new_n_n562_ | new_n_n563_;
  assign new_n_n556_ = new_n_n843_ | new_n_n844_ | new_n_n850_;
  assign new_n_n552_ = new_n_n555_ | new_n_n554_ | new_n_n652_;
  assign new_n_n544_ = new_n_n846_ | new_n_n865_ | new_n_n866_;
  assign new_n_n532_ = new_n_n889_ | new_n_n885_;
  assign new_n_n525_ = new_n_n792_ | new_n_n793_ | new_n_n794_;
  assign new_n_n472_ = new_n_n480_ | new_n_n479_ | new_n_n478_;
  assign new_n_n464_ = new_n_n797_ | new_n_n800_ | new_n_n803_;
  assign new_n_n459_ = new_n_n386_ | new_n_n468_ | new_n_n467_;
  assign new_n_n438_ = new_n_n300_ | new_n_n445_ | new_n_n444_;
  assign new_n_n430_ = new_n_n778_ | new_n_n781_ | new_n_n782_;
  assign new_n_n378_ = new_n_n814_ | new_n_n819_ | new_n_n820_;
  assign new_n_n369_ = new_n_n383_ | new_n_n382_ | new_n_n381_;
  assign new_n_n344_ = new_n_n805_ | new_n_n808_ | new_n_n810_;
  assign new_n_n335_ = new_n_n340_ | new_n_n650_ | new_n_n955_;
  assign new_n_n285_ = new_n_n290_ | new_n_n289_ | new_n_n288_;
  assign new_n_n277_ = new_n_n932_ | new_n_n928_;
  assign new_n_n761_ = new_n_n261_ & new_n_n260_ & new_n_n753_;
  assign new_n_n239_ = new_ni_23__ & new_n_n750_ & new_n_n747_;
  assign new_n_n790_ = new_n_n242_ & new_n_n228_ & new_n_n232_;
  assign new_n_n224_ = new_ni_21__ & new_ni_28__ & new_n_n747_;
  assign new_n_n824_ = new_n_n197_ & new_n_n199_ & new_n_n198_;
  assign new_n_n194_ = new_ni_21__ & new_ni_23__ & new_n_n750_;
  assign new_n_n181_ = new_n_n743_ & new_ni_18__ & new_ni_19__;
  assign new_n_n176_ = new_n_n743_ & new_n_n754_ & new_ni_19__;
  assign new_n_n145_ = new_n_n751_ & new_ni_28__ & new_n_n747_;
  assign new_n_n140_ = new_ni_5__ & new_n_n743_ & new_n_n752_;
  assign new_n_n887_ = new_n_n134_ & new_n_n218_ & new_n_n232_;
  assign new_n_n888_ = new_n_n129_ & new_n_n258_ & new_n_n214_;
  assign new_n_n124_ = new_ni_3__ & new_n_n732_ & new_n_n754_;
  assign new_n_n912_ = new_n_n89_ & new_n_n88_ & new_n_n208_;
  assign new_n_n916_ = new_n_n107_ & new_n_n215_ & new_n_n214_;
  assign new_n_n921_ = new_n_n76_ & new_n_n161_ & new_n_n75_;
  assign new_n_n924_ = new_n_n71_ & new_n_n161_ & new_n_n70_;
  assign new_no_42__ = 1'b0;
  assign new_n_n745_ = ~new_ni_11__;
  assign new_n_n738_ = ~new_ni_8__;
  assign new_n_n727_ = ~new_ni_15__;
  assign new_n_n720_ = ~new_ni_39__;
  assign new_n_n710_ = new_n_n759_ | new_n_n760_ | new_n_n761_;
  assign new_n_n660_ = new_n_n877_ | new_n_n879_ | new_n_n880_;
  assign new_n_n649_ = new_n_n949_ | new_n_n953_ | new_n_n954_;
  assign new_n_n642_ = new_n_n677_ | new_n_n676_ | new_n_n675_;
  assign new_n_n631_ = new_n_n646_ | new_n_n645_ | new_n_n644_;
  assign new_no_37__ = new_n_n625_ | new_n_n626_;
  assign new_n_n614_ = new_n_n907_ | new_n_n908_ | new_n_n909_;
  assign new_n_n564_ = new_n_n571_ | new_n_n570_ | new_n_n569_;
  assign new_no_30__ = new_n_n557_ | new_n_n558_;
  assign new_no_29__ = new_n_n553_ | new_n_n552_ | new_n_n277_;
  assign new_n_n541_ = new_n_n954_ | new_n_n931_;
  assign new_n_n535_ = new_n_n837_ | new_n_n838_ | new_n_n849_;
  assign new_n_n526_ = new_n_n786_ | new_n_n787_ | new_n_n790_;
  assign new_n_n475_ = new_n_n650_ | new_n_n489_ | new_n_n488_;
  assign new_n_n465_ = new_n_n787_ | new_n_n789_ | new_n_n790_;
  assign new_n_n458_ = new_n_n466_ | new_n_n465_ | new_n_n347_;
  assign new_n_n448_ = new_n_n785_ | new_n_n787_ | new_n_n790_;
  assign new_n_n431_ = new_n_n775_ | new_n_n776_ | new_n_n777_;
  assign new_n_n381_ = new_n_n795_ | new_n_n797_ | new_n_n802_;
  assign new_n_n370_ = new_n_n386_ | new_n_n385_ | new_n_n384_;
  assign new_no_15__ = new_n_n365_ | new_n_n364_ | new_n_n371_;
  assign new_n_n353_ = new_n_n356_ | new_n_n355_ | new_n_n354_;
  assign new_n_n288_ = new_n_n909_ | new_n_n920_ | new_no_41__;
  assign new_n_n278_ = new_n_n906_ | new_n_n907_ | new_n_n909_;
  assign new_n_n757_ = new_n_n70_ & new_n_n266_;
  assign new_n_n783_ = new_n_n236_ & new_n_n235_ & new_n_n234_;
  assign new_n_n229_ = new_n_n751_ & new_ni_26__ & new_ni_28__;
  assign new_n_n795_ = new_n_n268_ & new_n_n225_ & new_n_n240_;
  assign new_n_n189_ = new_ni_20__ & new_ni_21__ & new_ni_26__;
  assign new_n_n840_ = new_n_n183_ & new_n_n215_ & new_n_n214_;
  assign new_n_n845_ = new_n_n246_ & new_n_n177_ & new_n_n753_;
  assign new_n_n144_ = new_n_n146_ & new_n_n246_ & new_n_n145_;
  assign new_n_n880_ = new_n_n135_ & new_n_n178_ & new_n_n214_;
  assign new_n_n886_ = new_n_n169_ & new_n_n168_ & new_n_n130_;
  assign new_n_n913_ = new_n_n120_ & new_n_n148_ & new_n_n234_;
  assign new_n_n917_ = new_ni_30__ & new_n_n81_;
  assign new_n_n920_ = new_n_n78_ & new_n_n258_ & new_n_n77_;
  assign new_n_n70_ = new_ni_22__ & new_ni_29__ & new_n_n753_;
  assign new_no_43__ = new_no_44__ | new_n_n777_;
  assign new_n_n746_ = ~new_ni_27__;
  assign new_n_n737_ = ~new_ni_7__;
  assign new_n_n728_ = ~new_ni_1__;
  assign new_n_n719_ = ~new_ni_32__;
  assign new_n_n711_ = new_n_n755_ | new_n_n756_ | new_n_n757_;
  assign new_n_n659_ = new_n_n882_ | new_n_n885_ | new_n_n888_;
  assign new_n_n650_ = new_n_n941_ | new_n_n943_ | new_n_n944_;
  assign new_n_n641_ = new_n_n325_ | new_n_n674_ | new_n_n673_;
  assign new_n_n632_ = new_n_n486_ | new_n_n648_ | new_n_n647_;
  assign new_n_n624_ = new_n_n762_ | new_n_n764_ | new_n_n783_;
  assign new_n_n615_ = new_n_n900_ | new_n_n901_ | new_n_n903_;
  assign new_n_n563_ = new_n_n567_ | new_n_n566_ | new_n_n565_;
  assign new_n_n557_ = new_n_n909_ | new_n_n907_;
  assign new_n_n551_ = new_n_n765_ | new_n_n770_ | new_n_n771_;
  assign new_n_n542_ = new_n_n894_ | new_n_n904_ | new_n_n930_;
  assign new_n_n534_ = new_n_n851_ | new_n_n857_ | new_n_n858_;
  assign new_n_n527_ = new_n_n780_ | new_no_44__ | new_n_n782_;
  assign new_n_n474_ = new_n_n486_ | new_n_n485_ | new_n_n484_;
  assign new_n_n466_ = new_n_n783_ | new_n_n785_ | new_n_n786_;
  assign new_n_n457_ = new_n_n464_ | new_n_n463_ | new_n_n462_;
  assign new_n_n449_ = new_n_n779_ | new_n_n780_ | new_n_n783_;
  assign new_n_n440_ = new_n_n451_ | new_n_n450_ | new_n_n449_;
  assign new_n_n380_ = new_n_n803_ | new_n_n804_ | new_n_n805_;
  assign new_n_n371_ = new_n_n953_ | new_n_n952_;
  assign new_n_n363_ = new_n_n771_ | new_n_n772_ | new_n_n776_;
  assign new_n_n354_ = new_n_n576_ | new_n_n358_ | new_n_n357_;
  assign new_n_n287_ = new_n_n935_ | new_n_n938_ | new_n_n942_;
  assign new_n_n279_ = new_n_n898_ | new_n_n899_ | new_n_n903_;
  assign new_n_n272_ = new_n_n829_ | new_n_n835_ | new_n_n854_;
  assign new_n_n789_ = new_n_n246_ & new_n_n230_ & new_ni_30__;
  assign new_no_21__ = new_n_n255_ & new_n_n229_ & new_n_n234_;
  assign new_n_n225_ = new_n_n751_ & new_n_n746_ & new_ni_28__;
  assign new_n_n836_ = new_n_n182_ & new_n_n189_ & new_n_n264_;
  assign new_n_n183_ = new_n_n740_ & new_n_n754_ & new_n_n752_;
  assign new_n_n182_ = new_n_n745_ & new_ni_18__ & new_n_n752_;
  assign new_n_n139_ = new_ni_0__ & new_ni_10__ & new_n_n754_;
  assign new_n_n134_ = new_n_n735_ & new_n_n754_ & new_n_n752_;
  assign new_n_n130_ = new_ni_32__ & new_n_n734_;
  assign new_n_n87_ = new_n_n733_ & new_ni_15__ & new_n_n754_;
  assign new_n_n81_ = new_n_n82_ & new_n_n161_ & new_n_n50_;
  assign new_n_n76_ = new_n_n735_ & new_ni_3__ & new_ni_18__;
  assign new_n_n71_ = new_n_n735_ & new_n_n733_ & new_n_n754_;
  assign new_n_n702_ = new_n_n873_ | new_n_n881_ | new_n_n883_;
  assign new_n_n691_ = new_n_n696_ | new_n_n695_ | new_n_n694_;
  assign new_n_n681_ = new_n_n795_ | new_n_n796_ | new_n_n797_;
  assign new_n_n670_ = new_n_n840_ | new_n_n841_ | new_n_n842_;
  assign new_n_n605_ = new_n_n608_ | new_n_n607_ | new_n_n949_;
  assign new_n_n595_ = new_n_n849_ | new_n_n850_ | new_n_n852_;
  assign new_n_n584_ = new_n_n281_ | new_n_n280_ | new_n_n592_;
  assign new_n_n574_ = new_n_n835_ | new_n_n836_ | new_n_n839_;
  assign new_n_n517_ = new_n_n520_ | new_n_n519_ | new_n_n518_;
  assign new_n_n507_ = new_n_n799_ | new_n_n800_ | new_n_n801_;
  assign new_n_n496_ = new_n_n841_ | new_n_n842_ | new_n_n846_;
  assign new_n_n485_ = new_n_n687_ | new_n_n352_ | new_n_n432_;
  assign new_n_n469_ = new_n_n487_ | new_n_n471_;
  assign new_n_n411_ = new_n_n416_ | new_n_n415_ | new_n_n414_;
  assign new_n_n401_ = new_n_n826_ | new_n_n833_ | new_n_n837_;
  assign new_n_n390_ = new_n_n399_ | new_n_n374_ | new_n_n398_;
  assign new_n_n375_ = new_n_n855_ | new_n_n856_ | new_n_n857_;
  assign new_n_n364_ = new_n_n368_ | new_n_n367_ | new_n_n366_;
  assign new_n_n307_ = new_n_n310_ | new_n_n311_;
  assign new_n_n297_ = new_n_n871_ | new_n_n897_ | new_n_n937_;
  assign new_n_n283_ = new_n_n843_ | new_n_n844_ | new_n_n853_;
  assign new_n_n273_ = new_n_n804_ | new_n_n832_ | new_n_n834_;
  assign new_n_n266_ = new_ni_19__ & new_ni_20__ & new_ni_21__;
  assign new_n_n784_ = new_n_n69_ & new_n_n260_ & new_ni_30__;
  assign new_n_n792_ = new_n_n242_ & new_n_n227_ & new_n_n232_;
  assign new_n_n222_ = new_ni_21__ & new_ni_26__ & new_ni_30__;
  assign new_n_n215_ = new_n_n749_ & new_ni_21__ & new_ni_22__;
  assign new_n_n810_ = new_n_n216_ & new_n_n91_ & new_n_n234_;
  assign new_n_n179_ = new_ni_0__ & new_n_n754_ & new_n_n752_;
  assign new_n_n848_ = new_n_n263_ & new_n_n174_ & new_ni_30__;
  assign new_n_n855_ = new_n_n170_ & new_n_n141_ & new_n_n753_;
  assign new_n_n859_ = new_n_n164_ & new_n_n163_ & new_n_n269_;
  assign new_n_n863_ = new_n_n157_ & new_n_n215_ & new_n_n156_;
  assign new_n_n889_ = new_ni_30__ & new_n_n127_;
  assign new_n_n121_ = new_ni_33__ & new_n_n734_;
  assign new_n_n114_ = new_n_n115_ & new_n_n161_ & new_n_n260_;
  assign new_n_n902_ = new_n_n107_ & new_n_n207_ & new_n_n234_;
  assign new_n_n906_ = new_ni_30__ & new_n_n100_;
  assign new_n_n92_ = new_ni_21__ & new_n_n746_ & new_n_n750_;
  assign new_n_n3_ = new_n_n5_ & new_n_n6_;
  assign new_n_n701_ = new_n_n884_ | new_n_n887_ | new_n_n891_;
  assign new_n_n692_ = new_n_n699_ | new_n_n698_ | new_n_n697_;
  assign new_n_n680_ = new_n_n798_ | new_n_n800_ | new_n_n801_;
  assign new_n_n671_ = new_n_n837_ | new_n_n838_ | new_n_n839_;
  assign new_no_36__ = new_n_n605_ | new_n_n606_;
  assign new_n_n596_ = new_n_n840_ | new_n_n843_ | new_n_n844_;
  assign new_n_n583_ = new_n_n554_ | new_n_n591_ | new_n_n590_;
  assign new_n_n575_ = new_n_n827_ | new_n_n829_ | new_n_n832_;
  assign new_no_25__ = new_n_n904_ | new_n_n517_;
  assign new_n_n508_ = new_n_n796_ | new_n_n797_ | new_n_n798_;
  assign new_n_n495_ = new_n_n849_ | new_n_n851_ | new_n_n856_;
  assign new_n_n486_ = new_n_n711_ | new_n_n689_ | new_n_n688_;
  assign new_n_n460_ = new_n_n886_ | new_n_n895_ | new_n_n948_;
  assign new_n_n421_ = new_n_n836_ | new_n_n841_ | new_n_n855_;
  assign new_n_n400_ = new_n_n838_ | new_n_n840_ | new_n_n849_;
  assign new_n_n391_ = new_n_n675_ | new_n_n401_ | new_n_n400_;
  assign new_n_n374_ = new_n_n858_ | new_n_n859_ | new_n_n860_;
  assign new_n_n365_ = new_n_n486_ | new_n_n370_ | new_n_n369_;
  assign new_n_n306_ = new_n_n486_ | new_n_n309_ | new_n_n308_;
  assign new_n_n298_ = new_n_n836_ | new_n_n840_ | new_n_n848_;
  assign new_n_n282_ = new_n_n860_ | new_n_n867_ | new_n_n868_;
  assign new_no_6__ = new_n_n276_ | new_n_n275_ | new_n_n274_;
  assign new_n_n260_ = new_ni_22__ & new_n_n750_ & new_ni_29__;
  assign new_n_n780_ = new_n_n265_ & new_n_n239_ & new_ni_30__;
  assign new_n_n226_ = new_n_n751_ & new_ni_25__ & new_ni_30__;
  assign new_n_n798_ = new_n_n242_ & new_n_n223_ & new_n_n240_;
  assign new_n_n214_ = new_n_n750_ & new_n_n747_ & new_ni_30__;
  assign new_n_n809_ = new_n_n138_ & new_n_n212_;
  assign new_n_n178_ = new_ni_20__ & new_ni_21__ & new_ni_22__;
  assign new_n_n174_ = new_ni_21__ & new_ni_26__ & new_ni_29__;
  assign new_n_n169_ = new_n_n754_ & new_n_n752_ & new_ni_21__;
  assign new_n_n163_ = new_ni_20__ & new_n_n751_ & new_n_n746_;
  assign new_n_n151_ = new_n_n741_ & new_n_n744_ & new_n_n754_;
  assign new_n_n126_ = new_ni_5__ & new_ni_10__ & new_ni_18__;
  assign new_n_n894_ = new_n_n123_ & new_n_n122_ & new_n_n214_;
  assign new_n_n899_ = new_n_n753_ & new_n_n114_;
  assign new_n_n107_ = new_n_n728_ & new_n_n754_ & new_ni_19__;
  assign new_n_n99_ = new_ni_0__ & new_n_n742_ & new_ni_18__;
  assign new_n_n93_ = new_n_n725_ & new_n_n724_ & new_n_n739_;
  assign new_n_n4_ = new_n_n8_ & new_n_n223_ & new_n_n7_;
  assign new_n_n700_ = new_n_n896_ | new_n_n902_ | new_n_n905_;
  assign new_no_38__ = new_n_n940_ | new_n_n690_;
  assign new_n_n683_ = new_n_n784_ | new_n_n785_ | new_n_n786_;
  assign new_n_n672_ = new_n_n834_ | new_n_n835_ | new_n_n836_;
  assign new_n_n656_ = new_n_n899_ | new_n_n900_ | new_n_n901_;
  assign new_n_n604_ = new_n_n762_ | new_n_n764_ | new_n_n766_;
  assign new_n_n593_ = new_n_n868_ | new_n_n869_ | new_n_n870_;
  assign new_n_n586_ = new_n_n675_ | new_n_n597_ | new_n_n596_;
  assign new_n_n576_ = new_n_n823_ | new_n_n824_ | new_n_n826_;
  assign new_n_n561_ = new_n_n766_ | new_n_n795_ | new_n_n849_;
  assign new_n_n554_ = new_n_n899_ | new_n_n903_ | new_n_n906_;
  assign new_n_n516_ = new_n_n774_ | new_n_n775_ | new_n_n776_;
  assign new_n_n505_ = new_n_n805_ | new_n_n806_ | new_n_n807_;
  assign new_n_n498_ = new_n_n831_ | new_n_n833_ | new_n_n836_;
  assign new_n_n487_ = new_n_n955_ | new_n_n954_;
  assign new_n_n471_ = new_n_n477_ | new_n_n476_ | new_n_n475_;
  assign new_n_n461_ = new_n_n827_ | new_n_n833_ | new_n_n870_;
  assign new_n_n420_ = new_n_n908_ | new_n_n949_ | new_n_n951_;
  assign new_n_n410_ = new_n_n759_ | new_n_n764_ | new_n_n767_;
  assign new_n_n392_ = new_n_n404_ | new_n_n403_ | new_n_n402_;
  assign new_n_n377_ = new_no_20__ | new_n_n827_ | new_n_n837_;
  assign new_n_n366_ = new_n_n374_ | new_n_n373_ | new_n_n372_;
  assign new_n_n326_ = new_n_n817_ | new_n_n821_ | new_no_20__;
  assign new_n_n316_ = new_n_n769_ | new_n_n771_ | new_n_n781_;
  assign new_n_n284_ = new_n_n286_ | new_n_n287_;
  assign new_n_n274_ = new_n_n277_ | new_n_n652_;
  assign new_n_n766_ = new_n_n268_ & new_n_n256_ & new_ni_30__;
  assign new_n_n775_ = new_n_n244_ & new_n_n255_;
  assign new_n_n791_ = new_n_n250_ & new_n_n229_ & new_n_n247_;
  assign new_n_n223_ = new_ni_21__ & new_ni_22__ & new_n_n750_;
  assign new_n_n814_ = new_n_n216_ & new_n_n207_ & new_n_n234_;
  assign new_n_n820_ = new_n_n268_ & new_n_n202_ & new_n_n234_;
  assign new_n_n180_ = new_n_n749_ & new_ni_21__ & new_ni_25__;
  assign new_n_n847_ = new_n_n263_ & new_n_n175_ & new_ni_30__;
  assign new_n_n168_ = new_ni_23__ & new_ni_29__ & new_n_n753_;
  assign new_n_n157_ = new_ni_9__ & new_n_n754_ & new_n_n752_;
  assign new_n_n868_ = new_n_n179_ & new_n_n80_ & new_n_n217_;
  assign new_n_n128_ = new_ni_0__ & new_n_n741_ & new_n_n744_;
  assign new_n_n122_ = new_ni_20__ & new_ni_21__ & new_n_n731_;
  assign new_n_n113_ = new_n_n739_ & new_ni_18__ & new_n_n752_;
  assign new_n_n105_ = new_n_n106_ & new_n_n246_ & new_n_n175_;
  assign new_n_n101_ = new_ni_0__ & new_n_n733_ & new_n_n727_;
  assign new_n_n909_ = new_n_n753_ & new_n_n94_;
  assign new_n_n5_ = new_n_n721_ & new_n_n713_ & new_n_n714_;
  assign new_n_n699_ = new_n_n909_ | new_n_n910_ | new_n_n913_;
  assign new_n_n690_ = new_n_n693_ | new_n_n692_ | new_n_n691_;
  assign new_n_n682_ = new_n_n787_ | new_n_n788_ | new_n_n789_;
  assign new_n_n673_ = new_n_n831_ | new_n_n832_ | new_n_n833_;
  assign new_n_n646_ = new_n_n684_ | new_n_n683_ | new_n_n682_;
  assign new_n_n603_ = new_n_n768_ | new_n_n774_ | new_n_n777_;
  assign new_n_n594_ = new_n_n853_ | new_n_n859_ | new_n_n867_;
  assign new_n_n585_ = new_n_n595_ | new_n_n594_ | new_n_n593_;
  assign new_n_n577_ = new_n_n801_ | new_n_n806_ | new_n_n813_;
  assign new_n_n560_ = new_n_n860_ | new_n_n859_;
  assign new_n_n555_ = new_n_n877_ | new_n_n879_ | new_n_n889_;
  assign new_n_n515_ = new_n_n777_ | new_n_n778_ | new_n_n779_;
  assign new_n_n506_ = new_n_n802_ | new_n_n803_ | new_n_n804_;
  assign new_n_n497_ = new_n_n837_ | new_n_n838_ | new_n_n840_;
  assign new_n_n488_ = new_n_n951_ | new_n_n952_ | new_n_n953_;
  assign new_n_n470_ = new_n_n474_ | new_n_n473_ | new_n_n472_;
  assign new_n_n462_ = new_n_n810_ | new_n_n819_ | new_n_n820_;
  assign new_n_n419_ = new_n_n952_ | new_n_n953_ | new_n_n954_;
  assign new_no_17__ = new_n_n412_ | new_n_n411_ | new_n_n413_;
  assign new_n_n402_ = new_n_n819_ | new_n_n820_ | new_no_20__;
  assign new_n_n376_ = new_n_n838_ | new_n_n849_ | new_n_n851_;
  assign new_n_n367_ = new_n_n377_ | new_n_n376_ | new_n_n375_;
  assign new_n_n325_ = new_n_n825_ | new_n_n826_ | new_n_n827_;
  assign new_no_12__ = new_n_n317_ | new_n_n318_;
  assign new_no_8__ = new_n_n284_ | new_n_n285_;
  assign new_n_n275_ = new_n_n280_ | new_n_n279_ | new_n_n278_;
  assign new_n_n771_ = new_n_n251_ & new_n_n270_;
  assign new_n_n250_ = new_ni_18__ & new_ni_19__ & new_n_n749_;
  assign new_n_n227_ = new_n_n751_ & new_ni_22__ & new_n_n750_;
  assign new_n_n797_ = new_n_n268_ & new_n_n225_ & new_n_n247_;
  assign new_n_n206_ = new_ni_21__ & new_ni_22__ & new_ni_30__;
  assign new_n_n202_ = new_n_n751_ & new_ni_27__ & new_n_n750_;
  assign new_n_n842_ = new_n_n181_ & new_n_n180_ & new_ni_30__;
  assign new_n_n175_ = new_n_n751_ & new_n_n750_ & new_ni_29__;
  assign new_n_n162_ = new_ni_0__ & new_ni_3__ & new_ni_18__;
  assign new_n_n156_ = new_ni_30__ & new_n_n750_;
  assign new_n_n867_ = new_n_n152_ & new_n_n199_ & new_n_n269_;
  assign new_n_n127_ = new_n_n128_ & new_n_n263_ & new_n_n145_;
  assign new_n_n123_ = new_ni_5__ & new_ni_18__ & new_n_n752_;
  assign new_n_n112_ = new_n_n749_ & new_n_n751_ & new_n_n746_;
  assign new_n_n106_ = new_ni_0__ & new_n_n744_ & new_n_n733_;
  assign new_n_n100_ = new_n_n101_ & new_n_n258_ & new_n_n86_;
  assign new_n_n94_ = new_n_n96_ & new_n_n161_ & new_n_n95_;
  assign new_n_n6_ = new_n_n720_ & new_n_n715_ & new_n_n722_;
  assign new_n_n698_ = new_n_n916_ | new_n_n918_ | new_n_n919_;
  assign new_n_n688_ = new_n_n761_ | new_n_n762_ | new_n_n763_;
  assign new_n_n677_ = new_n_n817_ | new_n_n818_ | new_n_n819_;
  assign new_n_n666_ = new_n_n854_ | new_n_n857_ | new_n_n858_;
  assign new_n_n636_ = new_n_n660_ | new_n_n659_ | new_n_n658_;
  assign new_n_n602_ = new_n_n778_ | new_n_n779_ | new_n_n780_;
  assign new_n_n591_ = new_n_n907_ | new_n_n909_ | new_n_n915_;
  assign new_n_n580_ = new_n_n944_ | new_n_n583_;
  assign new_n_n570_ = new_n_n889_ | new_n_n897_ | new_n_n909_;
  assign new_n_n546_ = new_n_n825_ | new_n_n828_ | new_n_n830_;
  assign new_no_28__ = new_n_n537_ | new_n_n536_;
  assign new_n_n514_ = new_n_n780_ | new_no_44__ | new_n_n781_;
  assign new_n_n503_ = new_n_n811_ | new_n_n814_ | new_n_n816_;
  assign new_n_n492_ = new_n_n876_ | new_n_n885_ | new_n_n886_;
  assign new_n_n481_ = new_n_n507_ | new_n_n506_ | new_n_n505_;
  assign new_n_n453_ = new_n_n758_ | new_n_n760_ | new_n_n761_;
  assign new_n_n442_ = new_n_n948_ | new_n_n951_ | new_n_n952_;
  assign new_n_n432_ = new_n_n771_ | new_n_n772_ | new_n_n773_;
  assign new_n_n418_ = new_n_n434_ | new_n_n433_ | new_n_n432_;
  assign new_n_n408_ = new_n_n778_ | new_n_n779_ | new_no_44__;
  assign new_n_n397_ = new_n_n885_ | new_n_n889_ | new_n_n897_;
  assign new_no_16__ = new_n_n387_ | new_n_n388_;
  assign new_n_n358_ = new_n_n836_ | new_n_n848_ | new_n_n897_;
  assign new_n_n348_ = new_n_n787_ | new_no_21__ | new_n_n790_;
  assign new_n_n337_ = new_n_n346_ | new_n_n345_ | new_n_n344_;
  assign new_n_n327_ = new_n_n805_ | new_n_n810_ | new_n_n814_;
  assign new_n_n324_ = new_n_n830_ | new_n_n831_ | new_n_n836_;
  assign new_n_n314_ = new_n_n791_ | new_n_n797_ | new_n_n798_;
  assign new_n_n304_ = new_n_n772_ | new_n_n776_ | new_n_n778_;
  assign new_n_n293_ = new_n_n955_ | new_n_n650_;
  assign new_n_n755_ = new_n_n269_ & new_n_n270_;
  assign new_n_n262_ = new_ni_18__ & new_n_n752_ & new_n_n749_;
  assign new_n_n765_ = new_n_n252_ & new_n_n263_;
  assign new_n_n251_ = new_ni_28__ & new_ni_29__ & new_ni_30__;
  assign new_n_n249_ = new_n_n751_ & new_ni_22__ & new_ni_29__;
  assign new_n_n243_ = new_n_n751_ & new_ni_24__ & new_n_n747_;
  assign new_n_n781_ = new_n_n262_ & new_n_n238_ & new_ni_30__;
  assign new_n_n786_ = new_n_n250_ & new_n_n233_ & new_n_n232_;
  assign new_n_n218_ = new_ni_20__ & new_ni_21__ & new_ni_25__;
  assign new_n_n807_ = new_n_n263_ & new_n_n213_ & new_n_n753_;
  assign new_n_n813_ = new_n_n208_ & new_n_n265_;
  assign new_n_n819_ = new_n_n204_ & new_n_n203_ & new_n_n214_;
  assign new_n_n821_ = new_n_n149_ & new_n_n180_ & new_ni_30__;
  assign new_n_n826_ = new_n_n204_ & new_n_n203_ & new_n_n208_;
  assign new_n_n833_ = new_n_n193_ & new_n_n203_ & new_n_n214_;
  assign new_n_n186_ = new_n_n749_ & new_n_n751_ & new_n_n750_;
  assign new_n_n177_ = new_ni_21__ & new_ni_23__ & new_ni_29__;
  assign new_n_n853_ = new_n_n192_ & new_n_n207_ & new_n_n234_;
  assign new_n_n165_ = new_ni_3__ & new_ni_6__ & new_n_n754_;
  assign new_n_n158_ = new_n_n737_ & new_n_n736_ & new_ni_18__;
  assign new_n_n152_ = new_ni_0__ & new_n_n754_ & new_ni_19__;
  assign new_n_n872_ = new_ni_30__ & new_n_n144_;
  assign new_n_n877_ = new_n_n139_ & new_n_n258_ & new_n_n138_;
  assign new_n_n133_ = new_n_n749_ & new_ni_21__ & new_n_n750_;
  assign new_n_n125_ = new_n_n741_ & new_n_n732_ & new_n_n754_;
  assign new_n_n119_ = new_n_n750_ & new_ni_29__ & new_n_n730_;
  assign new_n_n117_ = new_ni_0__ & new_ni_10__ & new_ni_18__;
  assign new_n_n109_ = new_ni_20__ & new_n_n751_ & new_n_n729_;
  assign new_n_n904_ = new_ni_30__ & new_n_n102_;
  assign new_n_n95_ = new_n_n746_ & new_ni_28__ & new_ni_29__;
  assign new_n_n80_ = new_ni_20__ & new_n_n751_ & new_ni_23__;
  assign new_n_n922_ = new_n_n107_ & new_n_n74_ & new_n_n214_;
  assign new_n_n0_ = new_n_n2_ & new_n_n1_ & new_ni_44__;
  assign new_n_n697_ = new_n_n921_ | new_n_n922_ | new_n_n923_;
  assign new_n_n689_ = new_n_n758_ | new_n_n759_ | new_n_n760_;
  assign new_n_n676_ = new_n_n820_ | new_n_n821_ | new_no_20__;
  assign new_n_n667_ = new_n_n851_ | new_n_n852_ | new_n_n853_;
  assign new_n_n626_ = new_n_n632_ | new_n_n631_ | new_n_n630_;
  assign new_n_n601_ = new_n_n782_ | new_n_n783_ | new_n_n786_;
  assign new_n_n592_ = new_n_n892_ | new_n_n893_ | new_n_n898_;
  assign new_no_35__ = new_n_n582_ | new_n_n581_ | new_n_n580_;
  assign new_n_n571_ = new_n_n872_ | new_n_n874_ | new_n_n882_;
  assign new_n_n545_ = new_n_n831_ | new_n_n842_ | new_n_n845_;
  assign new_n_n536_ = new_n_n540_ | new_n_n539_ | new_n_n538_;
  assign new_n_n513_ = new_n_n782_ | new_n_n783_ | new_n_n784_;
  assign new_n_n504_ = new_n_n808_ | new_n_n809_ | new_n_n810_;
  assign new_n_n491_ = new_n_n889_ | new_n_n895_ | new_n_n897_;
  assign new_n_n482_ = new_n_n510_ | new_n_n509_ | new_n_n508_;
  assign new_n_n452_ = new_n_n762_ | new_n_n763_ | new_n_n766_;
  assign new_n_n443_ = new_n_n870_ | new_n_n878_ | new_n_n945_;
  assign new_n_n422_ = new_n_n824_ | new_n_n825_ | new_n_n826_;
  assign new_n_n417_ = new_n_n431_ | new_n_n430_ | new_n_n315_;
  assign new_n_n409_ = new_n_n772_ | new_n_n773_ | new_n_n776_;
  assign new_n_n396_ = new_n_n937_ | new_n_n941_ | new_n_n943_;
  assign new_n_n387_ = new_n_n391_ | new_n_n390_ | new_n_n389_;
  assign new_n_n357_ = new_n_n908_ | new_n_n937_ | new_n_n941_;
  assign new_n_n349_ = new_n_n779_ | new_n_n780_ | new_n_n786_;
  assign new_n_n336_ = new_n_n343_ | new_n_n342_ | new_n_n341_;
  assign new_n_n328_ = new_n_n799_ | new_n_n800_ | new_n_n802_;
  assign new_n_n323_ = new_n_n840_ | new_n_n841_ | new_n_n954_;
  assign new_n_n315_ = new_n_n783_ | new_n_n784_ | new_n_n785_;
  assign new_n_n303_ = new_n_n783_ | new_n_n785_ | new_no_21__;
  assign new_n_n294_ = new_n_n299_ | new_n_n298_ | new_n_n297_;
  assign new_n_n268_ = new_ni_18__ & new_ni_19__ & new_ni_20__;
  assign new_n_n759_ = new_n_n263_ & new_n_n174_ & new_n_n753_;
  assign new_n_n256_ = new_n_n751_ & new_ni_27__ & new_n_n747_;
  assign new_n_n770_ = new_n_n252_ & new_n_n268_;
  assign new_n_n772_ = new_n_n250_ & new_n_n249_ & new_ni_30__;
  assign new_n_n776_ = new_n_n250_ & new_n_n29_ & new_ni_30__;
  assign new_n_n237_ = new_ni_21__ & new_ni_23__ & new_n_n747_;
  assign new_n_n232_ = new_ni_30__ & new_n_n747_;
  assign new_n_n217_ = new_n_n750_ & new_ni_29__ & new_n_n753_;
  assign new_n_n213_ = new_n_n751_ & new_ni_24__ & new_ni_29__;
  assign new_n_n207_ = new_n_n749_ & new_n_n751_ & new_ni_22__;
  assign new_n_n203_ = new_ni_20__ & new_n_n751_ & new_ni_26__;
  assign new_no_20__ = new_n_n193_ & new_n_n203_ & new_n_n264_;
  assign new_n_n825_ = new_n_n254_ & new_n_n223_ & new_n_n234_;
  assign new_n_n192_ = new_ni_0__ & new_ni_18__ & new_ni_19__;
  assign new_n_n187_ = new_ni_3__ & new_n_n754_ & new_n_n752_;
  assign new_n_n172_ = new_ni_20__ & new_ni_21__ & new_ni_24__;
  assign new_n_n171_ = new_ni_10__ & new_n_n754_ & new_ni_19__;
  assign new_n_n857_ = new_n_n167_ & new_n_n166_ & new_n_n198_;
  assign new_n_n862_ = new_n_n158_ & new_n_n258_ & new_ni_28__;
  assign new_n_n866_ = new_n_n153_ & new_n_n258_ & new_ni_28__;
  assign new_n_n150_ = new_n_n752_ & new_n_n749_ & new_n_n751_;
  assign new_n_n137_ = new_ni_10__ & new_ni_18__ & new_n_n752_;
  assign new_n_n883_ = new_n_n134_ & new_n_n189_ & new_n_n232_;
  assign new_n_n892_ = new_n_n125_ & new_n_n166_ & new_n_n198_;
  assign new_n_n896_ = new_n_n120_ & new_n_n172_ & new_n_n232_;
  assign new_n_n116_ = new_ni_25__ & new_ni_29__ & new_n_n753_;
  assign new_n_n110_ = new_n_n739_ & new_n_n754_ & new_n_n752_;
  assign new_n_n905_ = new_n_n120_ & new_n_n207_ & new_n_n234_;
  assign new_n_n96_ = new_n_n735_ & new_n_n726_ & new_ni_18__;
  assign new_n_n918_ = new_n_n134_ & new_n_n80_ & new_n_n217_;
  assign new_n_n74_ = new_n_n749_ & new_ni_21__ & new_ni_23__;
  assign new_n_n1_ = new_n_n722_ & new_n_n721_ & new_n_n713_;
  assign new_n_n696_ = new_n_n924_ | new_n_n925_ | new_n_n926_;
  assign new_n_n686_ = new_n_n770_ | new_n_n771_ | new_n_n772_;
  assign new_n_n679_ = new_n_n811_ | new_n_n812_ | new_n_n813_;
  assign new_n_n668_ = new_n_n846_ | new_n_n849_ | new_n_n850_;
  assign new_n_n617_ = new_n_n868_ | new_n_n875_ | new_n_n879_;
  assign new_n_n600_ = new_n_n787_ | new_n_n792_ | new_n_n794_;
  assign new_n_n589_ = new_n_n711_ | new_n_n710_ | new_n_n604_;
  assign new_n_n582_ = new_n_n589_ | new_n_n588_ | new_n_n587_;
  assign new_n_n572_ = new_n_n863_ | new_n_n867_ | new_n_n871_;
  assign new_n_n529_ = new_n_n767_ | new_n_n768_ | new_n_n774_;
  assign new_n_n518_ = new_n_n523_ | new_n_n522_ | new_n_n521_;
  assign new_n_n512_ = new_n_n785_ | new_n_n786_ | new_n_n787_;
  assign new_n_n501_ = new_n_n821_ | new_no_20__ | new_n_n822_;
  assign new_n_n494_ = new_n_n857_ | new_n_n858_ | new_n_n859_;
  assign new_n_n483_ = new_n_n513_ | new_n_n512_ | new_n_n511_;
  assign new_n_n451_ = new_n_n767_ | new_n_n768_ | new_n_n769_;
  assign new_n_n434_ = new_n_n765_ | new_n_n766_ | new_n_n767_;
  assign new_n_n423_ = new_no_20__ | new_n_n822_ | new_n_n823_;
  assign new_n_n416_ = new_n_n429_ | new_n_n428_ | new_n_n427_;
  assign new_n_n406_ = new_n_n791_ | new_n_n794_ | new_n_n795_;
  assign new_n_n399_ = new_n_n851_ | new_n_n855_ | new_n_n857_;
  assign new_n_n388_ = new_n_n394_ | new_n_n393_ | new_n_n392_;
  assign new_n_n356_ = new_n_n363_ | new_n_n362_ | new_n_n361_;
  assign new_n_n346_ = new_n_n795_ | new_n_n799_ | new_n_n800_;
  assign new_n_n339_ = new_n_n352_ | new_n_n351_ | new_n_n350_;
  assign new_n_n329_ = new_n_n795_ | new_n_n797_ | new_n_n798_;
  assign new_n_n322_ = new_n_n687_ | new_n_n332_ | new_n_n304_;
  assign new_n_n312_ = new_n_n817_ | new_n_n825_ | new_n_n826_;
  assign new_no_11__ = new_n_n307_ | new_n_n306_;
  assign new_n_n295_ = new_n_n302_ | new_n_n301_ | new_n_n300_;
  assign new_n_n281_ = new_n_n872_ | new_n_n874_ | new_n_n877_;
  assign new_n_n267_ = new_ni_21__ & new_ni_29__ & new_n_n753_;
  assign new_n_n261_ = new_ni_18__ & new_ni_20__ & new_ni_21__;
  assign new_n_n257_ = new_ni_26__ & new_n_n750_ & new_ni_29__;
  assign new_n_n252_ = new_ni_21__ & new_ni_29__ & new_ni_30__;
  assign new_n_n248_ = new_ni_14__ & new_n_n746_ & new_n_n750_;
  assign new_n_n242_ = new_n_n754_ & new_ni_19__ & new_ni_20__;
  assign new_no_44__ = new_n_n263_ & new_n_n253_ & new_ni_30__;
  assign new_n_n785_ = new_n_n250_ & new_n_n233_ & new_n_n240_;
  assign new_n_n793_ = new_n_n226_ & new_n_n262_;
  assign new_n_n221_ = new_n_n744_ & new_ni_18__ & new_ni_19__;
  assign new_n_n802_ = new_n_n219_ & new_n_n218_ & new_n_n217_;
  assign new_n_n212_ = new_ni_18__ & new_n_n749_ & new_n_n751_;
  assign new_n_n812_ = new_n_n209_ & new_n_n210_;
  assign new_n_n204_ = new_ni_17__ & new_ni_18__ & new_n_n752_;
  assign new_n_n201_ = new_n_n751_ & new_n_n746_ & new_n_n750_;
  assign new_n_n196_ = new_n_n751_ & new_ni_26__ & new_n_n747_;
  assign new_n_n832_ = new_n_n152_ & new_n_n224_ & new_ni_30__;
  assign new_n_n837_ = new_n_n188_ & new_n_n186_ & new_n_n234_;
  assign new_n_n843_ = new_n_n179_ & new_n_n178_ & new_n_n232_;
  assign new_n_n849_ = new_n_n173_ & new_n_n163_ & new_n_n264_;
  assign new_n_n854_ = new_n_n171_ & new_n_n235_ & new_n_n232_;
  assign new_n_n164_ = new_ni_4__ & new_ni_18__ & new_ni_19__;
  assign new_n_n159_ = new_n_n738_ & new_ni_16__ & new_ni_18__;
  assign new_n_n153_ = new_ni_7__ & new_n_n736_ & new_ni_18__;
  assign new_n_n869_ = new_n_n151_ & new_n_n150_ & new_n_n232_;
  assign new_n_n143_ = new_ni_0__ & new_ni_18__ & new_n_n752_;
  assign new_n_n882_ = new_n_n192_ & new_n_n136_ & new_n_n198_;
  assign new_n_n890_ = new_n_n126_ & new_n_n258_ & new_n_n214_;
  assign new_n_n120_ = new_n_n735_ & new_ni_18__ & new_ni_19__;
  assign new_n_n898_ = new_n_n117_ & new_n_n37_ & new_n_n116_;
  assign new_n_n901_ = new_n_n110_ & new_n_n109_ & new_n_n108_;
  assign new_n_n103_ = new_ni_25__ & new_n_n750_ & new_n_n747_;
  assign new_n_n908_ = new_ni_33__ & new_n_n97_;
  assign new_no_32__ = new_n_n93_ & new_n_n92_ & new_n_n247_;
  assign new_n_n85_ = new_n_n87_ & new_n_n266_ & new_n_n86_;
  assign new_n_n2_ = new_n_n730_ & new_n_n720_ & new_n_n715_;
  assign new_n_n695_ = new_n_n927_ | new_n_n929_ | new_n_n933_;
  assign new_n_n687_ = new_n_n764_ | new_n_n765_ | new_n_n766_;
  assign new_n_n678_ = new_n_n814_ | new_n_n815_ | new_n_n816_;
  assign new_n_n669_ = new_n_n843_ | new_n_n844_ | new_n_n845_;
  assign new_n_n607_ = new_n_n614_ | new_n_n613_ | new_n_n612_;
  assign new_n_n599_ = new_n_n800_ | new_n_n802_ | new_n_n803_;
  assign new_n_n590_ = new_no_41__ | new_n_n928_ | new_n_n932_;
  assign new_n_n581_ = new_n_n586_ | new_n_n585_ | new_n_n584_;
  assign new_n_n573_ = new_n_n841_ | new_n_n852_ | new_n_n854_;
  assign new_n_n528_ = new_n_n775_ | new_n_n777_ | new_n_n779_;
  assign new_n_n519_ = new_n_n526_ | new_n_n525_ | new_n_n524_;
  assign new_n_n511_ = new_n_n788_ | new_n_n789_ | new_no_21__;
  assign new_n_n502_ = new_n_n817_ | new_n_n819_ | new_n_n820_;
  assign new_n_n493_ = new_n_n860_ | new_n_n871_ | new_n_n872_;
  assign new_n_n484_ = new_n_n516_ | new_n_n515_ | new_n_n514_;
  assign new_n_n441_ = new_n_n711_ | new_n_n453_ | new_n_n452_;
  assign new_n_n433_ = new_n_n768_ | new_n_n769_ | new_n_n770_;
  assign new_n_n424_ = new_n_n819_ | new_n_n820_ | new_n_n821_;
  assign new_n_n415_ = new_n_n426_ | new_n_n425_ | new_n_n424_;
  assign new_n_n407_ = new_n_n786_ | new_no_21__ | new_n_n790_;
  assign new_n_n398_ = new_n_n870_ | new_n_n871_ | new_n_n872_;
  assign new_n_n389_ = new_n_n397_ | new_n_n396_ | new_n_n395_;
  assign new_n_n355_ = new_n_n360_ | new_n_n344_ | new_n_n359_;
  assign new_n_n347_ = new_n_n791_ | new_n_n792_ | new_n_n794_;
  assign new_n_n338_ = new_n_n349_ | new_n_n348_ | new_n_n347_;
  assign new_n_n330_ = new_n_n785_ | new_no_21__ | new_n_n791_;
  assign new_n_n321_ = new_n_n331_ | new_n_n330_ | new_n_n329_;
  assign new_n_n313_ = new_n_n800_ | new_n_n803_ | new_n_n808_;
  assign new_n_n305_ = new_n_n764_ | new_n_n766_ | new_n_n769_;
  assign new_n_n296_ = new_n_n305_ | new_n_n304_ | new_n_n303_;
  assign new_no_5__ = new_n_n850_ | new_n_n273_;
  assign new_n_n756_ = new_n_n267_ & new_n_n268_;
  assign new_n_n760_ = new_n_n262_ & new_n_n238_ & new_n_n753_;
  assign new_n_n764_ = new_n_n258_ & new_n_n257_ & new_n_n753_;
  assign new_n_n769_ = new_n_n269_ & new_n_n265_;
  assign new_n_n247_ = new_n_n753_ & new_n_n747_;
  assign new_n_n777_ = new_n_n263_ & new_n_n243_ & new_ni_30__;
  assign new_n_n238_ = new_ni_21__ & new_n_n750_ & new_ni_29__;
  assign new_n_n233_ = new_n_n751_ & new_ni_26__ & new_n_n750_;
  assign new_n_n794_ = new_n_n268_ & new_n_n201_ & new_n_n232_;
  assign new_n_n799_ = new_n_n222_ & new_n_n250_;
  assign new_n_n216_ = new_ni_1__ & new_n_n754_ & new_ni_19__;
  assign new_n_n808_ = new_n_n216_ & new_n_n74_ & new_n_n214_;
  assign new_n_n208_ = new_ni_28__ & new_n_n747_ & new_n_n753_;
  assign new_n_n818_ = new_n_n205_ & new_n_n262_;
  assign new_n_n822_ = new_n_n268_ & new_n_n201_ & new_n_n234_;
  assign new_n_n827_ = new_n_n204_ & new_n_n203_ & new_n_n217_;
  assign new_n_n193_ = new_n_n742_ & new_ni_18__ & new_n_n752_;
  assign new_n_n188_ = new_ni_5__ & new_n_n754_ & new_n_n752_;
  assign new_n_n844_ = new_n_n179_ & new_n_n189_ & new_n_n232_;
  assign new_n_n173_ = new_ni_5__ & new_ni_18__ & new_ni_19__;
  assign new_n_n170_ = new_ni_13__ & new_n_n739_ & new_ni_21__;
  assign new_n_n858_ = new_n_n165_ & new_n_n166_ & new_n_n198_;
  assign new_n_n861_ = new_n_n159_ & new_n_n258_ & new_ni_28__;
  assign new_n_n865_ = new_n_n154_ & new_n_n258_ & new_ni_28__;
  assign new_n_n149_ = new_ni_10__ & new_ni_18__ & new_ni_19__;
  assign new_n_n873_ = new_n_n73_ & new_n_n224_ & new_ni_30__;
  assign new_n_n138_ = new_ni_25__ & new_n_n747_ & new_ni_30__;
  assign new_n_n891_ = new_n_n134_ & new_n_n172_ & new_n_n232_;
  assign new_n_n895_ = new_n_n169_ & new_n_n168_ & new_n_n121_;
  assign new_n_n115_ = new_ni_0__ & new_n_n733_ & new_n_n754_;
  assign new_n_n108_ = new_n_n746_ & new_n_n747_ & new_n_n753_;
  assign new_n_n102_ = new_n_n104_ & new_n_n258_ & new_n_n103_;
  assign new_n_n97_ = new_n_n157_ & new_n_n215_ & new_n_n214_;
  assign new_n_n91_ = new_n_n749_ & new_n_n751_ & new_ni_23__;
  assign new_n_n86_ = new_ni_22__ & new_n_n750_ & new_n_n747_;
  assign new_n_n954_ = new_n_n3_ & new_n_n4_;
  assign new_n_n928_ = new_n_n753_ & new_n_n67_;
  assign new_n_n59_ = new_n_n17_ & new_n_n26_ & new_n_n235_;
  assign new_n_n935_ = new_ni_30__ & new_n_n52_;
  assign new_n_n938_ = new_ni_30__ & new_n_n44_;
  assign new_n_n36_ = new_n_n38_ & new_n_n37_ & new_n_n57_;
  assign new_n_n67_ = new_n_n68_ & new_n_n166_ & new_n_n257_;
  assign new_n_n932_ = new_n_n232_ & new_n_n59_;
  assign new_n_n52_ = new_n_n53_ & new_n_n166_ & new_n_n57_;
  assign new_n_n43_ = new_n_n735_ & new_n_n744_ & new_n_n733_;
  assign new_n_n37_ = new_ni_19__ & new_n_n749_ & new_n_n751_;
  assign new_n_n68_ = new_ni_0__ & new_ni_17__ & new_ni_18__;
  assign new_n_n58_ = new_n_n735_ & new_ni_11__ & new_ni_18__;
  assign new_n_n50_ = new_n_n746_ & new_n_n750_ & new_ni_29__;
  assign new_n_n45_ = new_ni_21__ & new_ni_25__ & new_n_n747_;
  assign new_n_n38_ = new_ni_0__ & new_n_n745_ & new_ni_18__;
  assign new_n_n927_ = new_n_n66_ & new_n_n69_ & new_n_n214_;
  assign new_n_n57_ = new_ni_26__ & new_ni_28__ & new_n_n747_;
  assign new_n_n51_ = new_n_n735_ & new_n_n733_ & new_ni_18__;
  assign new_n_n44_ = new_n_n30_ & new_n_n263_ & new_n_n45_;
  assign new_n_n941_ = new_n_n39_ & new_n_n118_;
  assign new_n_n955_ = new_n_n0_ & new_n_n19_;
  assign new_n_n685_ = new_n_n773_ | new_n_n774_ | new_n_n775_;
  assign new_n_n674_ = new_n_n828_ | new_n_n829_ | new_n_n830_;
  assign new_n_n578_ = new_n_n781_ | new_n_n784_ | new_n_n785_;
  assign new_n_n69_ = new_ni_18__ & new_n_n752_ & new_ni_21__;
  assign new_n_n32_ = new_n_n753_ & new_n_n734_ & new_n_n719_;
  assign new_n_n947_ = new_n_n232_ & new_n_n24_;
  assign new_n_n15_ = new_n_n17_ & new_n_n16_ & new_n_n218_;
  assign new_n_n8_ = new_n_n740_ & new_n_n754_ & new_n_n749_;
  assign new_n_n684_ = new_n_n781_ | new_n_n782_ | new_n_n783_;
  assign new_n_n675_ = new_n_n822_ | new_n_n823_ | new_n_n824_;
  assign new_n_n587_ = new_n_n600_ | new_n_n599_ | new_n_n598_;
  assign new_n_n926_ = new_n_n120_ & new_n_n136_ & new_n_n217_;
  assign new_n_n31_ = new_ni_34__ & new_n_n723_;
  assign new_n_n24_ = new_n_n27_ & new_n_n26_ & new_n_n25_;
  assign new_n_n950_ = new_n_n214_ & new_n_n15_;
  assign new_n_n953_ = new_n_n9_ & new_n_n19_;
  assign new_n_n703_ = new_n_n706_ | new_n_n705_ | new_n_n885_;
  assign new_n_n693_ = new_n_n702_ | new_n_n701_ | new_n_n700_;
  assign new_n_n597_ = new_n_n832_ | new_n_n833_ | new_n_n834_;
  assign new_n_n945_ = new_n_n31_ & new_n_n22_;
  assign new_n_n22_ = new_n_n246_ & new_n_n177_ & new_n_n32_;
  assign new_n_n17_ = new_ni_0__ & new_n_n733_ & new_ni_10__;
  assign new_n_n9_ = new_n_n2_ & new_n_n10_ & new_n_n714_;
  assign new_no_39__ = new_n_n589_ | new_n_n704_ | new_n_n703_;
  assign new_n_n694_ = new_n_n934_ | new_n_n936_ | new_n_n939_;
  assign new_n_n606_ = new_n_n611_ | new_n_n610_ | new_n_n609_;
  assign new_n_n30_ = new_ni_0__ & new_ni_10__ & new_n_n745_;
  assign new_n_n23_ = new_n_n723_ & new_n_n718_ & new_ni_35__;
  assign new_n_n16_ = new_n_n745_ & new_n_n727_ & new_n_n752_;
  assign new_n_n10_ = new_n_n722_ & new_n_n721_ & new_ni_43__;
  assign new_n_n722_ = ~new_ni_41__;
  assign new_no_40__ = new_n_n535_ | new_n_n712_ | new_n_n894_;
  assign new_n_n616_ = new_n_n888_ | new_n_n898_ | new_n_n899_;
  assign new_n_n49_ = new_n_n51_ & new_n_n161_ & new_n_n50_;
  assign new_n_n939_ = new_n_n753_ & new_n_n42_;
  assign new_n_n943_ = new_n_n35_ & new_n_n118_;
  assign new_n_n27_ = new_ni_0__ & new_n_n733_ & new_n_n745_;
  assign new_n_n18_ = new_n_n20_ & new_n_n21_;
  assign new_n_n952_ = new_n_n11_ & new_n_n22_;
  assign new_n_n721_ = ~new_ni_42__;
  assign new_n_n712_ = new_n_n851_ | new_n_n880_ | new_n_n890_;
  assign new_n_n625_ = new_n_n629_ | new_n_n628_ | new_n_n627_;
  assign new_n_n936_ = new_ni_30__ & new_n_n49_;
  assign new_n_n42_ = new_n_n43_ & new_n_n246_ & new_n_n175_;
  assign new_n_n34_ = new_n_n730_ & new_ni_39__ & new_n_n722_;
  assign new_n_n946_ = new_n_n753_ & new_n_n28_;
  assign new_n_n949_ = new_n_n18_ & new_n_n19_;
  assign new_n_n11_ = new_n_n12_ & new_n_n13_;
  assign new_n_n742_ = ~new_ni_17__;
  assign new_n_n731_ = ~new_ni_25__;
  assign new_n_n635_ = new_n_n657_ | new_n_n656_ | new_n_n655_;
  assign new_n_n63_ = new_ni_8__ & new_ni_16__ & new_n_n754_;
  assign new_n_n933_ = new_ni_30__ & new_n_n56_;
  assign new_n_n33_ = new_ni_42__ & new_n_n34_;
  assign new_n_n25_ = new_ni_21__ & new_ni_26__ & new_n_n750_;
  assign new_n_n20_ = new_n_n721_ & new_n_n722_;
  assign new_n_n12_ = new_ni_37__ & new_n_n716_;
  assign new_n_n741_ = ~new_ni_2__;
  assign new_n_n732_ = ~new_ni_6__;
  assign new_n_n645_ = new_n_n428_ | new_n_n525_ | new_n_n681_;
  assign new_n_n62_ = new_n_n63_ & new_n_n266_ & new_n_n184_;
  assign new_n_n56_ = new_n_n58_ & new_n_n166_ & new_n_n57_;
  assign new_n_n944_ = new_n_n33_ & new_n_n19_;
  assign new_n_n26_ = new_n_n727_ & new_n_n752_ & new_ni_20__;
  assign new_n_n19_ = new_n_n183_ & new_n_n215_ & new_n_n217_;
  assign new_n_n13_ = new_n_n723_ & new_n_n718_ & new_n_n717_;
  assign new_n_n751_ = ~new_ni_21__;
  assign new_n_n655_ = new_n_n903_ | new_n_n904_ | new_n_n906_;
  assign new_n_n929_ = new_n_n66_ & new_n_n65_ & new_n_n64_;
  assign new_n_n930_ = new_n_n753_ & new_n_n62_;
  assign new_n_n54_ = new_n_n55_ & new_n_n263_ & new_n_n145_;
  assign new_n_n46_ = new_n_n157_ & new_n_n215_ & new_n_n48_;
  assign new_n_n39_ = new_ni_39__ & new_n_n722_ & new_n_n721_;
  assign new_n_n948_ = new_n_n23_ & new_n_n22_;
  assign new_n_n951_ = new_n_n14_ & new_n_n22_;
  assign new_no_1__ = new_n_n896_ | new_n_n891_;
  assign new_n_n752_ = ~new_ni_19__;
  assign new_n_n665_ = new_n_n859_ | new_n_n860_ | new_n_n861_;
  assign new_n_n64_ = new_ni_22__ & new_n_n747_ & new_ni_30__;
  assign new_n_n61_ = new_ni_7__ & new_n_n736_ & new_n_n754_;
  assign new_n_n55_ = new_n_n735_ & new_ni_2__ & new_n_n744_;
  assign new_n_n937_ = new_n_n47_ & new_n_n46_;
  assign new_n_n940_ = new_ni_30__ & new_n_n40_;
  assign new_n_n21_ = new_n_n730_ & new_n_n720_ & new_ni_40__;
  assign new_n_n14_ = new_ni_36__ & new_n_n13_;
  assign new_n_n65_ = new_n_n754_ & new_ni_20__ & new_ni_21__;
  assign new_n_n60_ = new_n_n61_ & new_n_n266_ & new_n_n184_;
  assign new_n_n53_ = new_ni_0__ & new_ni_11__ & new_ni_18__;
  assign new_n_n48_ = new_n_n750_ & new_ni_30__ & new_n_n734_;
  assign new_n_n40_ = new_n_n41_ & new_n_n246_ & new_n_n145_;
  assign new_n_n942_ = new_ni_30__ & new_n_n36_;
  assign new_n_n28_ = new_n_n30_ & new_n_n250_ & new_n_n29_;
  assign new_n_n66_ = new_n_n735_ & new_n_n733_ & new_n_n727_;
  assign new_n_n931_ = new_n_n753_ & new_n_n60_;
  assign new_n_n934_ = new_ni_30__ & new_n_n54_;
  assign new_n_n47_ = new_ni_39__ & new_n_n723_;
  assign new_n_n41_ = new_n_n735_ & new_n_n741_ & new_n_n744_;
  assign new_n_n35_ = new_n_n720_ & new_n_n722_ & new_ni_42__;
  assign new_n_n29_ = new_n_n751_ & new_ni_25__ & new_ni_29__;
endmodule


