// Benchmark "adder10" written by ABC on Sat Apr 29 10:28:08 2023

module adder10 ( 
    a9, a8, a7, a6, a5, a4, a3, a2, a1, a0, b9, b8, b7, b6, b5, b4, b3, b2,
    b1, b0, cin,
    cout, s9, s8, s7, s6, s5, s4, s3, s2, s1, s0  );
  input  a9, a8, a7, a6, a5, a4, a3, a2, a1, a0, b9, b8, b7, b6, b5, b4,
    b3, b2, b1, b0, cin;
  output cout, s9, s8, s7, s6, s5, s4, s3, s2, s1, s0;
  assign cout = (((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2) & (b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6) & (a7 | b7) & (a8 | b8) & (b9 | a9)) | ((b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6) & (a7 | b7) & (a8 | b8) & (b9 | a9) & ((a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | ((b5 | a5) & (a6 | b6) & (a7 | b7) & (a8 | b8) & (b9 | a9) & ((a4 & (b4 | (b3 & a3))) | (b3 & a3 & b4))) | ((a7 | b7) & (a8 | b8) & (b9 | a9) & ((a6 & (b6 | (b5 & a5))) | (b5 & a5 & b6))) | ((b9 | a9) & ((a8 & (b8 | (a7 & b7))) | (a7 & b7 & b8))) | (b9 & a9);
  assign s9 = ((~b9 ^ a9) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2) & (b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6) & (a7 | b7) & (a8 | b8)) | ((b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6) & (a7 | b7) & (a8 | b8) & ((a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | ((b5 | a5) & (a6 | b6) & (a7 | b7) & (a8 | b8) & ((a4 & (b4 | (b3 & a3))) | (b3 & a3 & b4))) | ((a7 | b7) & (a8 | b8) & ((a6 & (b6 | (b5 & a5))) | (b5 & a5 & b6))) | (a8 & (b8 | (a7 & b7))) | (a7 & b7 & b8))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (b9 ^ a9) & (~b1 | ~a1) & (~a2 | ~b2) & (~b3 | ~a3) & (~a4 | ~b4) & (~b5 | ~a5) & (~a6 | ~b6) & (~a7 | ~b7) & (~a8 | ~b8)) | (((~a2 & (~b2 | (~b1 & ~a1))) | (~b1 & ~a1 & ~b2)) & (b9 ^ a9) & (~b3 | ~a3) & (~a4 | ~b4) & (~b5 | ~a5) & (~a6 | ~b6) & (~a7 | ~b7) & (~a8 | ~b8)) | (((~a4 & (~b4 | (~b3 & ~a3))) | (~b3 & ~a3 & ~b4)) & (b9 ^ a9) & (~b5 | ~a5) & (~a6 | ~b6) & (~a7 | ~b7) & (~a8 | ~b8)) | (((~a6 & (~b6 | (~b5 & ~a5))) | (~b5 & ~a5 & ~b6)) & (b9 ^ a9) & (~a7 | ~b7) & (~a8 | ~b8)) | ((b9 ^ a9) & ((~a8 & (~b8 | (~a7 & ~b7))) | (~a7 & ~b7 & ~b8)));
  assign s8 = ((~a8 ^ b8) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2) & (b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6) & (a7 | b7)) | ((b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6) & (a7 | b7) & ((a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | ((b5 | a5) & (a6 | b6) & (a7 | b7) & ((a4 & (b4 | (b3 & a3))) | (b3 & a3 & b4))) | ((a7 | b7) & ((a6 & (b6 | (b5 & a5))) | (b5 & a5 & b6))) | (a7 & b7))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (a8 ^ b8) & (~b1 | ~a1) & (~a2 | ~b2) & (~b3 | ~a3) & (~a4 | ~b4) & (~b5 | ~a5) & (~a7 | ~b7) & (~a6 | ~b6)) | (((~a2 & (~b2 | (~b1 & ~a1))) | (~b1 & ~a1 & ~b2)) & (a8 ^ b8) & (~b3 | ~a3) & (~a4 | ~b4) & (~b5 | ~a5) & (~a7 | ~b7) & (~a6 | ~b6)) | (((~a4 & (~b4 | (~b3 & ~a3))) | (~b3 & ~a3 & ~b4)) & (a8 ^ b8) & (~b5 | ~a5) & (~a7 | ~b7) & (~a6 | ~b6)) | (((~a6 & (~b6 | (~b5 & ~a5))) | (~b5 & ~a5 & ~b6)) & (~a7 | ~b7) & (a8 ^ b8)) | (~a7 & ~b7 & (a8 ^ b8));
  assign s7 = ((~a7 ^ b7) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2) & (b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6)) | ((b3 | a3) & (a4 | b4) & (b5 | a5) & (a6 | b6) & ((a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | ((b5 | a5) & (a6 | b6) & ((a4 & (b4 | (b3 & a3))) | (b3 & a3 & b4))) | (a6 & (b6 | (b5 & a5))) | (b5 & a5 & b6))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (a7 ^ b7) & (~b1 | ~a1) & (~a2 | ~b2) & (~b3 | ~a3) & (~a4 | ~b4) & (~b5 | ~a5) & (~a6 | ~b6)) | (((~a2 & (~b2 | (~b1 & ~a1))) | (~b1 & ~a1 & ~b2)) & (a7 ^ b7) & (~b3 | ~a3) & (~a4 | ~b4) & (~b5 | ~a5) & (~a6 | ~b6)) | (((~a4 & (~b4 | (~b3 & ~a3))) | (~b3 & ~a3 & ~b4)) & (a7 ^ b7) & (~b5 | ~a5) & (~a6 | ~b6)) | ((a7 ^ b7) & ((~a6 & (~b6 | (~b5 & ~a5))) | (~b5 & ~a5 & ~b6)));
  assign s6 = ((~a6 ^ b6) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2) & (b3 | a3) & (a4 | b4) & (b5 | a5)) | ((b3 | a3) & (a4 | b4) & (b5 | a5) & ((a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | ((b5 | a5) & ((a4 & (b4 | (b3 & a3))) | (b3 & a3 & b4))) | (b5 & a5))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (a6 ^ b6) & (~b1 | ~a1) & (~a2 | ~b2) & (~b3 | ~a3) & (~b5 | ~a5) & (~a4 | ~b4)) | (((~a2 & (~b2 | (~b1 & ~a1))) | (~b1 & ~a1 & ~b2)) & (a6 ^ b6) & (~b3 | ~a3) & (~b5 | ~a5) & (~a4 | ~b4)) | (((~a4 & (~b4 | (~b3 & ~a3))) | (~b3 & ~a3 & ~b4)) & (~b5 | ~a5) & (a6 ^ b6)) | (~b5 & ~a5 & (a6 ^ b6));
  assign s5 = ((~b5 ^ a5) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2) & (b3 | a3) & (a4 | b4)) | ((b3 | a3) & (a4 | b4) & ((a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | (a4 & (b4 | (b3 & a3))) | (b3 & a3 & b4))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (b5 ^ a5) & (~b1 | ~a1) & (~a2 | ~b2) & (~b3 | ~a3) & (~a4 | ~b4)) | (((~a2 & (~b2 | (~b1 & ~a1))) | (~b1 & ~a1 & ~b2)) & (b5 ^ a5) & (~b3 | ~a3) & (~a4 | ~b4)) | ((b5 ^ a5) & ((~a4 & (~b4 | (~b3 & ~a3))) | (~b3 & ~a3 & ~b4)));
  assign s4 = ((a4 ^ ~b4) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2) & (b3 | a3)) | ((b3 | a3) & ((a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | (b3 & a3))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (a4 ^ b4) & (~b1 | ~a1) & (~b3 | ~a3) & (~a2 | ~b2)) | (((~a2 & (~b2 | (~b1 & ~a1))) | (~b1 & ~a1 & ~b2)) & (~b3 | ~a3) & (a4 ^ b4)) | (~b3 & ~a3 & (a4 ^ b4));
  assign s3 = ((b3 ^ ~a3) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1) & (a2 | b2)) | (a2 & (b2 | (b1 & a1))) | (b1 & a1 & b2))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (b3 ^ a3) & (~b1 | ~a1) & (~a2 | ~b2)) | ((b3 ^ a3) & ((~a2 & (~b2 | (~b1 & ~a1))) | (~b1 & ~a1 & ~b2)));
  assign s2 = ((a2 ^ ~b2) & ((((cin & (a0 | b0)) | (a0 & b0)) & (b1 | a1)) | (b1 & a1))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (~b1 | ~a1) & (a2 ^ b2)) | (~b1 & ~a1 & (a2 ^ b2));
  assign s1 = ((b1 ^ ~a1) & ((cin & (a0 | b0)) | (a0 & b0))) | (((~a0 & ~b0) | (~cin & (~a0 | ~b0))) & (b1 ^ a1));
  assign s0 = cin ? (a0 ^ ~b0) : (a0 ^ b0);
endmodule


