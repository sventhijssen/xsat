// Benchmark "top" written by ABC on Fri Mar 31 12:13:24 2023

module top ( 
    pa1, pb2, pc3, pd4, pe5, pp, pa0, pb3, pc2, pd5, pe4, pq, pa3, pb0,
    pc1, pf4, pg5, pr, pa2, pb1, pc0, pf5, pg4, ps, pa5, pd0, pe1, pf2,
    pg3, pt, pa4, pd1, pe0, pf3, pg2, pu, pb4, pc5, pd2, pe3, pf0, pg1, pv,
    pb5, pc4, pd3, pe2, pf1, pg0, pw, ph0, pi1, pj2, pk3, pl4, pm5, ph1,
    pi0, pj3, pk2, pl5, pm4, py, ph2, pi3, pj0, pk1, pn4, po5, pz, ph3,
    pi2, pj1, pk0, pn5, po4, ph4, pi5, pl0, pm1, pn2, po3, ph5, pi4, pl1,
    pm0, pn3, po2, pj4, pk5, pl2, pm3, pn0, po1, pj5, pk4, pl3, pm2, pn1,
    po0, pp0, pq1, pr2, ps3, pt4, pa, pp1, pq0, pr3, ps2, pu4, pb, pp2,
    pq3, pr0, ps1, pv4, pc, pp3, pq2, pr1, ps0, pw4, pd, pp4, pq5, pt0,
    pu1, pv2, pw3, pe, pp5, pq4, pt1, pu0, pv3, pw2, pf, pr4, pt2, pu3,
    pv0, pw1, pg, pr5, ps4, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1,
    py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, px4, pm, py4, pn,
    pz4, po,
    pf6, pg7, ph8, pi9, pq10, pf7, pg6, ph9, pi8, pp10, pd6, pe7, pj8, pk9,
    ps10, pd7, pe6, pj9, pk8, pr10, pb6, pc7, pl8, pm9, pu10, pb7, pc6,
    pl9, pm8, pt10, pa7, pn8, po9, pw10, pa6, pn9, po8, pv10, pa9, pn6,
    po7, py10, pa8, pn7, po6, px10, pb8, pc9, pl6, pm7, pb9, pc8, pl7, pm6,
    pd8, pe9, pj6, pk7, pd9, pe8, pj7, pk6, pf8, pg9, ph6, pi7, pf9, pg8,
    ph7, pi6, pa10, pu5, pv6, pw7, px8, py9, pt5, pv7, pw6, px9, py8, pc10,
    pt6, pu7, pw5, pz8, pb10, pt7, pu6, pv5, pz9, pe10, pr6, ps7, pd10,
    pr7, ps6, pg10, pp6, pq7, ps5, pf10, pp7, pq6, pi10, pp8, pq9, ph10,
    pp9, pq8, pk10, pr8, ps9, pj10, pr9, ps8, pm10, pt8, pu9, py5, pz6,
    pl10, pt9, pu8, px5, pz7, po10, pv8, pw9, px6, py7, pn10, pv9, pw8,
    px7, py6, pz5  );
  input  pa1, pb2, pc3, pd4, pe5, pp, pa0, pb3, pc2, pd5, pe4, pq, pa3,
    pb0, pc1, pf4, pg5, pr, pa2, pb1, pc0, pf5, pg4, ps, pa5, pd0, pe1,
    pf2, pg3, pt, pa4, pd1, pe0, pf3, pg2, pu, pb4, pc5, pd2, pe3, pf0,
    pg1, pv, pb5, pc4, pd3, pe2, pf1, pg0, pw, ph0, pi1, pj2, pk3, pl4,
    pm5, ph1, pi0, pj3, pk2, pl5, pm4, py, ph2, pi3, pj0, pk1, pn4, po5,
    pz, ph3, pi2, pj1, pk0, pn5, po4, ph4, pi5, pl0, pm1, pn2, po3, ph5,
    pi4, pl1, pm0, pn3, po2, pj4, pk5, pl2, pm3, pn0, po1, pj5, pk4, pl3,
    pm2, pn1, po0, pp0, pq1, pr2, ps3, pt4, pa, pp1, pq0, pr3, ps2, pu4,
    pb, pp2, pq3, pr0, ps1, pv4, pc, pp3, pq2, pr1, ps0, pw4, pd, pp4, pq5,
    pt0, pu1, pv2, pw3, pe, pp5, pq4, pt1, pu0, pv3, pw2, pf, pr4, pt2,
    pu3, pv0, pw1, pg, pr5, ps4, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi,
    px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, px4, pm, py4,
    pn, pz4, po;
  output pf6, pg7, ph8, pi9, pq10, pf7, pg6, ph9, pi8, pp10, pd6, pe7, pj8,
    pk9, ps10, pd7, pe6, pj9, pk8, pr10, pb6, pc7, pl8, pm9, pu10, pb7,
    pc6, pl9, pm8, pt10, pa7, pn8, po9, pw10, pa6, pn9, po8, pv10, pa9,
    pn6, po7, py10, pa8, pn7, po6, px10, pb8, pc9, pl6, pm7, pb9, pc8, pl7,
    pm6, pd8, pe9, pj6, pk7, pd9, pe8, pj7, pk6, pf8, pg9, ph6, pi7, pf9,
    pg8, ph7, pi6, pa10, pu5, pv6, pw7, px8, py9, pt5, pv7, pw6, px9, py8,
    pc10, pt6, pu7, pw5, pz8, pb10, pt7, pu6, pv5, pz9, pe10, pr6, ps7,
    pd10, pr7, ps6, pg10, pp6, pq7, ps5, pf10, pp7, pq6, pi10, pp8, pq9,
    ph10, pp9, pq8, pk10, pr8, ps9, pj10, pr9, ps8, pm10, pt8, pu9, py5,
    pz6, pl10, pt9, pu8, px5, pz7, po10, pv8, pw9, px6, py7, pn10, pv9,
    pw8, px7, py6, pz5;
  wire new_na1_, new_nb2_, new_nc3_, new_nd4_, new_ne5_, new_np_, new_na0_,
    new_nb3_, new_nc2_, new_nd5_, new_ne4_, new_nq_, new_na3_, new_nb0_,
    new_nc1_, new_nf4_, new_ng5_, new_nr_, new_na2_, new_nb1_, new_nc0_,
    new_nf5_, new_ng4_, new_ns_, new_na5_, new_nd0_, new_ne1_, new_nf2_,
    new_ng3_, new_nt_, new_na4_, new_nd1_, new_ne0_, new_nf3_, new_ng2_,
    new_nu_, new_nb4_, new_nc5_, new_nd2_, new_ne3_, new_nf0_, new_ng1_,
    new_nv_, new_nb5_, new_nc4_, new_nd3_, new_ne2_, new_nf1_, new_ng0_,
    new_nw_, new_nh0_, new_ni1_, new_nj2_, new_nk3_, new_nl4_, new_nm5_,
    new_nh1_, new_ni0_, new_nj3_, new_nk2_, new_nl5_, new_nm4_, new_ny_,
    new_nh2_, new_ni3_, new_nj0_, new_nk1_, new_nn4_, new_no5_, new_nz_,
    new_nh3_, new_ni2_, new_nj1_, new_nk0_, new_nn5_, new_no4_, new_nh4_,
    new_ni5_, new_nl0_, new_nm1_, new_nn2_, new_no3_, new_nh5_, new_ni4_,
    new_nl1_, new_nm0_, new_nn3_, new_no2_, new_nj4_, new_nk5_, new_nl2_,
    new_nm3_, new_nn0_, new_no1_, new_nj5_, new_nk4_, new_nl3_, new_nm2_,
    new_nn1_, new_no0_, new_np0_, new_nq1_, new_nr2_, new_ns3_, new_nt4_,
    new_na_, new_np1_, new_nq0_, new_nr3_, new_ns2_, new_nu4_, new_nb_,
    new_np2_, new_nq3_, new_nr0_, new_ns1_, new_nv4_, new_nc_, new_np3_,
    new_nq2_, new_nr1_, new_ns0_, new_nw4_, new_nd_, new_np4_, new_nq5_,
    new_nt0_, new_nu1_, new_nv2_, new_nw3_, new_ne_, new_np5_, new_nq4_,
    new_nt1_, new_nu0_, new_nv3_, new_nw2_, new_nf_, new_nr4_, new_nt2_,
    new_nu3_, new_nv0_, new_nw1_, new_ng_, new_nr5_, new_ns4_, new_nt3_,
    new_nu2_, new_nv1_, new_nw0_, new_nh_, new_nx0_, new_ny1_, new_nz2_,
    new_ni_, new_nx1_, new_ny0_, new_nz3_, new_nj_, new_nx2_, new_ny3_,
    new_nz0_, new_nk_, new_nx3_, new_ny2_, new_nz1_, new_nl_, new_nx4_,
    new_nm_, new_ny4_, new_nn_, new_nz4_, new_no_, new_nf7_, new_nq7_,
    new_ny7_, new_ng8_, new_n_n1384_, new_nz8_, new_nk9_, new_nv9_,
    new_nj17_, new_nt17_, new_ne18_, new_nw18_, new_nq19_, new_n_n1314_,
    new_nb35_, new_nm35_, new_n_n1071_, new_n_n1064_, new_n_n1060_,
    new_nn39_, new_n_n1047_, new_n_n1024_, new_n_n1017_, new_ne42_,
    new_n_n1005_, new_n_n998_, new_n_n991_, new_ne43_, new_nm43_,
    new_ni44_, new_nt44_, new_na45_, new_n_n942_, new_ns45_, new_ny45_,
    new_n_n920_, new_n_n912_, new_n_n909_, new_n_n890_, new_n_n884_,
    new_nv49_, new_n_n877_, new_nz50_, new_nl51_, new_nq51_, new_n_n859_,
    new_nj52_, new_n_n849_, new_n_n841_, new_no53_, new_nl54_, new_nw54_,
    new_nh55_, new_ns55_, new_nd56_, new_no56_, new_nz56_, new_n_n785_,
    new_n_n774_, new_n_n763_, new_n_n752_, new_n_n741_, new_n_n730_,
    new_n_n719_, new_n_n708_, new_n_n686_, new_n_n675_, new_n_n664_,
    new_n_n654_, new_n_n643_, new_n_n632_, new_n_n621_, new_n_n610_,
    new_n_n599_, new_n_n588_, new_n_n577_, new_n_n566_, new_n_n555_,
    new_n_n544_, new_n_n533_, new_n_n522_, new_n_n511_, new_n_n500_,
    new_n_n489_, new_n_n478_, new_n_n467_, new_n_n456_, new_n_n445_,
    new_n_n434_, new_n_n423_, new_n_n412_, new_n_n401_, new_n_n390_,
    new_n_n368_, new_n_n357_, new_n_n346_, new_n_n335_, new_n_n324_,
    new_n_n313_, new_n_n302_, new_n_n291_, new_n_n258_, new_n_n247_,
    new_n_n236_, new_n_n225_, new_n_n214_, new_n_n203_, new_n_n192_,
    new_n_n149_, new_n_n138_, new_n_n127_, new_n_n116_, new_n_n105_,
    new_n_n94_, new_nu6_, new_nr7_, new_nx7_, new_nh8_, new_nq8_, new_na9_,
    new_nj9_, new_nw9_, new_nl17_, new_n_n1367_, new_n_n1360_, new_nu18_,
    new_nu19_, new_n_n1322_, new_nc35_, new_nl35_, new_nq38_, new_n_n1065_,
    new_n_n1059_, new_n_n1054_, new_nk40_, new_n_n1023_, new_nx41_,
    new_ng42_, new_n_n1006_, new_n_n997_, new_nx42_, new_ng43_,
    new_n_n979_, new_nv43_, new_nv44_, new_n_n948_, new_no45_, new_n_n935_,
    new_nb46_, new_n_n921_, new_np46_, new_nx46_, new_ns48_, new_n_n885_,
    new_n_n883_, new_n_n878_, new_na51_, new_nk51_, new_n_n867_, new_nv51_,
    new_nk52_, new_n_n850_, new_n_n840_, new_nn53_, new_nm54_, new_nv54_,
    new_ni55_, new_nr55_, new_ne56_, new_nn56_, new_n_n808_, new_n_n784_,
    new_n_n775_, new_n_n762_, new_n_n753_, new_n_n740_, new_n_n731_,
    new_n_n718_, new_n_n709_, new_n_n685_, new_n_n676_, new_n_n663_,
    new_nv10_, new_n_n642_, new_n_n633_, new_n_n620_, new_n_n611_,
    new_n_n589_, new_n_n587_, new_n_n578_, new_n_n565_, new_n_n556_,
    new_n_n543_, new_n_n534_, new_n_n521_, new_n_n512_, new_n_n499_,
    new_n_n490_, new_n_n488_, new_n_n466_, new_n_n457_, new_n_n444_,
    new_n_n435_, new_n_n422_, new_n_n413_, new_n_n400_, new_n_n391_,
    new_n_n367_, new_n_n358_, new_n_n345_, new_n_n336_, new_n_n323_,
    new_n_n314_, new_n_n301_, new_n_n292_, new_n_n268_, new_n_n246_,
    new_n_n237_, new_n_n224_, new_n_n215_, new_n_n202_, new_n_n193_,
    new_n_n148_, new_n_n139_, new_n_n126_, new_n_n117_, new_n_n104_,
    new_n_n95_, new_nf6_, new_nh6_, new_ns7_, new_na8_, new_ne8_, new_np8_,
    new_nb9_, new_nm9_, new_nt9_, new_no16_, new_n_n1375_, new_n_n1359_,
    new_ny18_, new_nm19_, new_nn22_, new_n_n1129_, new_nz34_, new_nk35_,
    new_n_n1073_, new_nu38_, new_nh39_, new_nt39_, new_nj40_, new_n_n1025_,
    new_nv41_, new_nh42_, new_n_n1004_, new_ns42_, new_nv42_, new_nq43_,
    new_n_n965_, new_n_n954_, new_n_n946_, new_nk45_, new_n_n936_,
    new_nd46_, new_n_n919_, new_n_n914_, new_n_n910_, new_n_n899_,
    new_n_n896_, new_n_n882_, new_nf50_, new_nv50_, new_nj51_, new_n_n869_,
    new_nu51_, new_nl52_, new_nv52_, new_n_n843_, new_nm53_, new_nj54_,
    new_nu54_, new_nj55_, new_nu55_, new_nb56_, new_nm56_, new_n_n798_,
    new_n_n787_, new_n_n776_, new_n_n761_, new_n_n750_, new_n_n743_,
    new_n_n732_, new_n_n699_, new_n_n688_, new_n_n677_, new_n_n662_,
    new_n_n652_, new_n_n645_, new_n_n634_, new_n_n619_, new_n_n601_,
    new_n_n590_, new_n_n564_, new_n_n553_, new_n_n546_, new_n_n535_,
    new_n_n520_, new_n_n509_, new_n_n502_, new_n_n491_, new_n_n465_,
    new_n_n454_, new_n_n447_, new_n_n436_, new_n_n421_, new_n_n410_,
    new_n_n403_, new_n_n392_, new_n_n366_, new_n_n355_, new_n_n348_,
    new_n_n337_, new_n_n322_, new_n_n311_, new_n_n304_, new_n_n293_,
    new_n_n267_, new_n_n256_, new_n_n238_, new_n_n223_, new_n_n212_,
    new_n_n205_, new_n_n194_, new_n_n169_, new_n_n158_, new_n_n125_,
    new_n_n114_, new_n_n107_, new_n_n96_, new_ng6_, new_nt7_, new_nz7_,
    new_nf8_, new_no8_, new_nc9_, new_nl9_, new_nu9_, new_nq16_,
    new_n_n1376_, new_nj18_, new_nx18_, new_no19_, new_nb22_, new_ny31_,
    new_na35_, new_nj35_, new_n_n1072_, new_n_n1066_, new_n_n1053_,
    new_n_n1048_, new_ni40_, new_ns41_, new_n_n1018_, new_nj42_, new_no42_,
    new_n_n999_, new_n_n992_, new_n_n972_, new_n_n966_, new_n_n953_,
    new_n_n947_, new_nn45_, new_nr45_, new_n_n926_, new_nh46_, new_n_n913_,
    new_n_n911_, new_n_n898_, new_n_n897_, new_nx49_, new_n_n876_,
    new_ny50_, new_ni51_, new_n_n868_, new_n_n860_, new_nm52_, new_n_n848_,
    new_n_n842_, new_nk53_, new_nk54_, new_nt54_, new_nk55_, new_nt55_,
    new_nc56_, new_nl56_, new_n_n788_, new_n_n786_, new_n_n777_,
    new_n_n760_, new_n_n751_, new_n_n742_, new_n_n733_, new_n_n698_,
    new_n_n689_, new_n_n687_, new_n_n661_, new_n_n653_, new_n_n644_,
    new_n_n635_, new_n_n609_, new_n_n600_, new_n_n591_, new_n_n563_,
    new_n_n554_, new_n_n545_, new_n_n536_, new_n_n519_, new_n_n510_,
    new_n_n501_, new_n_n492_, new_n_n464_, new_n_n455_, new_n_n446_,
    new_n_n437_, new_n_n420_, new_n_n411_, new_n_n402_, new_n_n393_,
    new_n_n365_, new_n_n356_, new_n_n347_, new_n_n338_, new_n_n321_,
    new_n_n312_, new_n_n303_, new_n_n294_, new_n_n266_, new_n_n257_,
    new_n_n248_, new_n_n222_, new_n_n213_, new_n_n204_, new_n_n195_,
    new_n_n168_, new_n_n159_, new_n_n124_, new_n_n115_, new_n_n106_,
    new_n_n97_, new_nd6_, new_nu7_, new_n_n1387_, new_nk8_, new_ns8_,
    new_nv8_, new_ng9_, new_nr9_, new_nr16_, new_n_n1374_, new_n_n1371_,
    new_ny17_, new_ni19_, new_nt21_, new_n_n1131_, new_n_n1124_, new_nx34_,
    new_ni35_, new_nn38_, new_n_n1067_, new_nn40_, new_nv40_, new_n_n1030_,
    new_nk42_, new_np42_, new_n_n986_, new_n_n981_, new_n_n974_,
    new_n_n967_, new_nw44_, new_ne45_, new_np45_, new_nu45_, new_nv45_,
    new_n_n923_, new_n_n915_, new_nw46_, new_ny47_, new_n_n895_,
    new_n_n888_, new_nm49_, new_nr50_, new_ng51_, new_n_n864_, new_n_n857_,
    new_ne52_, new_nt52_, new_n_n845_, new_ni53_, new_np54_, new_na55_,
    new_nd55_, new_no55_, new_nz55_, new_nk56_, new_n_n781_, new_n_n770_,
    new_n_n767_, new_n_n756_, new_n_n745_, new_n_n734_, new_n_n682_,
    new_n_n671_, new_n_n657_, new_n_n647_, new_n_n636_, new_n_n584_,
    new_n_n573_, new_n_n548_, new_n_n537_, new_n_n485_, new_n_n474_,
    new_n_n438_, new_n_n419_, new_n_n386_, new_n_n375_, new_n_n320_,
    new_n_n309_, new_n_n287_, new_n_n276_, new_n_n221_, new_n_n210_,
    new_n_n199_, new_n_n188_, new_n_n177_, new_n_n123_, new_n_n112_,
    new_n_n101_, new_n_n90_, new_nb6_, new_ne6_, new_nv7_, new_nb8_,
    new_nl8_, new_nr8_, new_nw8_, new_nf9_, new_ns9_, new_nl16_, new_nz16_,
    new_no17_, new_nv17_, new_nk19_, new_no21_, new_n_n1130_, new_n_n1125_,
    new_ny34_, new_nh35_, new_np38_, new_n_n1068_, new_np40_, new_nt40_,
    new_nr41_, new_n_n1009_, new_n_n1003_, new_n_n985_, new_n_n982_,
    new_n_n973_, new_nu43_, new_n_n952_, new_n_n945_, new_n_n939_,
    new_n_n932_, new_n_n929_, new_n_n924_, new_nk46_, new_nv46_, new_na48_,
    new_nl48_, new_ny48_, new_nj49_, new_nt50_, new_nf51_, new_n_n863_,
    new_nz51_, new_nf52_, new_n_n852_, new_n_n844_, new_nh53_, new_nq54_,
    new_nz54_, new_ne55_, new_nn55_, new_na56_, new_nj56_, new_n_n780_,
    new_n_n771_, new_n_n766_, new_n_n757_, new_n_n744_, new_n_n735_,
    new_n_n681_, new_n_n672_, new_n_n667_, new_n_n646_, new_n_n637_,
    new_n_n583_, new_n_n574_, new_n_n547_, new_n_n538_, new_n_n484_,
    new_n_n475_, new_n_n448_, new_n_n409_, new_n_n385_, new_n_n376_,
    new_n_n319_, new_n_n310_, new_n_n286_, new_n_n277_, new_n_n220_,
    new_n_n211_, new_n_n189_, new_n_n187_, new_n_n178_, new_n_n122_,
    new_n_n113_, new_n_n100_, new_n_n91_, new_nw7_, new_n_n1385_, new_ni8_,
    new_n_n1382_, new_nx8_, new_ni9_, new_np9_, new_n_n1379_, new_nb17_,
    new_nm17_, new_n_n1365_, new_n_n1362_, new_ns18_, new_nb21_,
    new_n_n1178_, new_nv28_, new_np31_, new_n_n1126_, new_nv34_, new_ng35_,
    new_nt38_, new_n_n1041_, new_nc41_, new_n_n1026_, new_nt42_,
    new_n_n989_, new_n_n984_, new_n_n980_, new_np43_, new_ns43_,
    new_n_n951_, new_n_n943_, new_n_n941_, new_n_n933_, new_n_n928_,
    new_ng46_, new_nj46_, new_nu46_, new_nb48_, new_no48_, new_nv48_,
    new_ni49_, new_nt49_, new_nc50_, new_n_n866_, new_nw51_, new_n_n855_,
    new_n_n851_, new_n_n846_, new_ng53_, new_nn54_, new_ny54_, new_nf55_,
    new_nq55_, new_nx55_, new_ni56_, new_n_n783_, new_n_n772_, new_n_n765_,
    new_n_n754_, new_n_n747_, new_n_n736_, new_n_n684_, new_n_n673_,
    new_n_n666_, new_n_n655_, new_n_n638_, new_n_n586_, new_n_n575_,
    new_n_n568_, new_n_n557_, new_n_n487_, new_n_n476_, new_n_n458_,
    new_n_n399_, new_n_n388_, new_n_n377_, new_n_n300_, new_n_n289_,
    new_n_n278_, new_n_n219_, new_n_n201_, new_n_n190_, new_n_n121_,
    new_n_n110_, new_n_n103_, new_n_n92_, new_nc6_, new_n_n1390_,
    new_n_n1386_, new_nj8_, new_n_n1383_, new_ny8_, new_nh9_, new_nq9_,
    new_ns16_, new_n_n1373_, new_n_n1372_, new_n_n1366_, new_n_n1361_,
    new_nr18_, new_n_n1345_, new_n_n1177_, new_n_n1175_, new_nr31_,
    new_nx31_, new_nw34_, new_nf35_, new_n_n1074_, new_n_n1036_,
    new_n_n1031_, new_np41_, new_n_n996_, new_n_n990_, new_na43_,
    new_nl43_, new_n_n975_, new_n_n968_, new_n_n950_, new_n_n944_,
    new_n_n940_, new_n_n934_, new_n_n927_, new_n_n922_, new_n_n916_,
    new_nt46_, new_nc48_, new_n_n894_, new_n_n889_, new_ng49_, new_nu49_,
    new_n_n879_, new_n_n865_, new_n_n858_, new_ni52_, new_nu52_, new_ny52_,
    new_nf53_, new_no54_, new_nx54_, new_ng55_, new_np55_, new_ny55_,
    new_nh56_, new_n_n782_, new_n_n773_, new_n_n764_, new_n_n755_,
    new_n_n746_, new_n_n737_, new_n_n683_, new_n_n674_, new_n_n665_,
    new_n_n656_, new_n_n648_, new_n_n585_, new_n_n576_, new_n_n567_,
    new_n_n558_, new_n_n486_, new_n_n477_, new_n_n468_, new_n_n389_,
    new_n_n387_, new_n_n378_, new_n_n299_, new_n_n290_, new_n_n288_,
    new_n_n209_, new_n_n200_, new_n_n191_, new_n_n120_, new_n_n111_,
    new_n_n102_, new_n_n93_, new_np6_, new_nc7_, new_nn7_, new_nb10_,
    new_no10_, new_ng16_, new_n_n1353_, new_nd29_, new_n_n1163_,
    new_n_n1121_, new_nr32_, new_ny32_, new_n_n1105_, new_no33_, new_np35_,
    new_na36_, new_n_n1099_, new_nz36_, new_n_n1088_, new_n_n1082_,
    new_nf38_, new_n_n1075_, new_n_n1058_, new_no39_, new_na40_,
    new_n_n1044_, new_n_n1037_, new_nx40_, new_no41_, new_ny42_, new_nj43_,
    new_n_n976_, new_n_n969_, new_ny43_, new_nn44_, new_ns46_, new_n_n905_,
    new_n_n902_, new_nr53_, new_n_n836_, new_ng54_, new_n_n817_, new_nr56_,
    new_nc57_, new_n_n804_, new_n_n793_, new_n_n727_, new_n_n716_,
    new_n_n705_, new_n_n694_, new_n_n678_, new_n_n618_, new_n_n607_,
    new_n_n596_, new_n_n580_, new_n_n569_, new_n_n508_, new_n_n497_,
    new_n_n481_, new_n_n470_, new_n_n459_, new_n_n398_, new_n_n382_,
    new_n_n371_, new_n_n360_, new_n_n349_, new_n_n283_, new_n_n272_,
    new_n_n261_, new_n_n250_, new_n_n239_, new_n_n184_, new_n_n174_,
    new_n_n163_, new_n_n152_, new_n_n141_, new_n_n130_, new_nx5_, new_no6_,
    new_nd7_, new_nm7_, new_no9_, new_na10_, new_nq10_, new_nf16_,
    new_n_n1356_, new_ne29_, new_nn29_, new_n_n1120_, new_nq32_,
    new_n_n1111_, new_n_n1106_, new_ny33_, new_nq35_, new_nz35_, new_no36_,
    new_ns36_, new_nh37_, new_nn37_, new_ng38_, new_nm38_, new_nb39_,
    new_nq39_, new_nw39_, new_nm40_, new_n_n1038_, new_nz40_, new_nm41_,
    new_n_n988_, new_nh43_, new_nn43_, new_n_n970_, new_ne44_, new_n_n955_,
    new_n_n917_, new_ng47_, new_n_n903_, new_ns53_, new_nc54_, new_n_n826_,
    new_n_n818_, new_ns56_, new_nb57_, new_n_n803_, new_n_n794_,
    new_n_n726_, new_n_n717_, new_n_n704_, new_n_n695_, new_n_n668_,
    new_n_n628_, new_n_n606_, new_n_n597_, new_n_n579_, new_n_n570_,
    new_n_n507_, new_n_n498_, new_n_n480_, new_n_n471_, new_n_n449_,
    new_n_n408_, new_n_n381_, new_n_n372_, new_n_n359_, new_n_n350_,
    new_n_n282_, new_n_n273_, new_n_n260_, new_n_n251_, new_n_n229_,
    new_n_n183_, new_n_n175_, new_n_n162_, new_n_n153_, new_n_n140_,
    new_n_n131_, new_ny5_, new_ns6_, new_na7_, new_nl7_, new_ne9_,
    new_nd10_, new_nm10_, new_nb16_, new_nt29_, new_n_n1151_, new_n_n1119_,
    new_nt32_, new_n_n1112_, new_ne33_, new_ni34_, new_nr35_, new_nc36_,
    new_n_n1100_, new_n_n1094_, new_nj37_, new_no37_, new_nd38_,
    new_n_n1076_, new_nc39_, new_ni39_, new_nu39_, new_n_n1043_, new_ns40_,
    new_n_n1033_, new_ng41_, new_n_n1020_, new_nz41_, new_n_n987_,
    new_n_n983_, new_n_n978_, new_nr43_, new_n_n961_, new_n_n956_,
    new_ne46_, new_nd47_, new_nr47_, new_nu53_, new_n_n834_, new_n_n828_,
    new_nh54_, new_nr54_, new_nt56_, new_ne57_, new_n_n806_, new_n_n795_,
    new_n_n779_, new_n_n768_, new_n_n725_, new_n_n714_, new_n_n707_,
    new_n_n696_, new_n_n680_, new_n_n669_, new_n_n627_, new_n_n616_,
    new_n_n598_, new_n_n582_, new_n_n571_, new_n_n528_, new_n_n517_,
    new_n_n483_, new_n_n472_, new_n_n439_, new_n_n418_, new_n_n384_,
    new_n_n373_, new_n_n340_, new_n_n329_, new_n_n285_, new_n_n274_,
    new_n_n259_, new_n_n241_, new_n_n230_, new_n_n186_, new_nv6_,
    new_n_n161_, new_n_n150_, new_n_n143_, new_n_n132_, new_nz5_, new_nq6_,
    new_nb7_, new_nk7_, new_nu8_, new_nc10_, new_nn10_, new_ny10_,
    new_nv29_, new_n_n1152_, new_ne32_, new_ns32_, new_nw32_, new_nc33_,
    new_ns34_, new_ns35_, new_nb36_, new_nn36_, new_n_n1095_, new_n_n1087_,
    new_n_n1081_, new_ne38_, new_n_n1077_, new_n_n1062_, new_n_n1057_,
    new_n_n1052_, new_n_n1042_, new_nr40_, new_n_n1032_, new_n_n1027_,
    new_n_n1019_, new_n_n1013_, new_nz42_, new_nk43_, new_n_n977_,
    new_n_n971_, new_n_n960_, new_nl44_, new_n_n930_, new_n_n906_,
    new_np47_, new_nv53_, new_n_n835_, new_n_n827_, new_n_n819_, new_nb55_,
    new_nu56_, new_nd57_, new_n_n805_, new_n_n796_, new_n_n778_,
    new_n_n769_, new_n_n724_, new_n_n715_, new_n_n706_, new_n_n697_,
    new_n_n679_, new_n_n670_, new_n_n626_, new_n_n617_, new_n_n608_,
    new_n_n581_, new_n_n572_, new_n_n527_, new_n_n518_, new_n_n482_,
    new_n_n473_, new_n_n429_, new_n_n428_, new_n_n383_, new_n_n374_,
    new_n_n339_, new_n_n330_, new_n_n284_, new_n_n275_, new_n_n249_,
    new_n_n240_, new_n_n231_, new_n_n185_, new_n_n176_, new_n_n160_,
    new_n_n151_, new_n_n142_, new_n_n133_, new_na6_, new_nj6_, new_ny6_,
    new_nj7_, new_nn8_, new_nk10_, new_nx10_, new_np30_, new_n_n1146_,
    new_n_n1118_, new_nk33_, new_nv33_, new_ng34_, new_nr34_, new_nt35_,
    new_ne36_, new_n_n1097_, new_ne37_, new_n_n1091_, new_n_n1084_,
    new_nt37_, new_n_n1078_, new_nr38_, new_nd39_, new_nm39_, new_n_n1050_,
    new_nh40_, new_n_n1040_, new_n_n1034_, new_n_n1028_, new_n_n1021_,
    new_n_n1014_, new_n_n1012_, new_n_n1008_, new_n_n1000_, new_n_n993_,
    new_nw43_, new_n_n957_, new_n_n937_, new_n_n907_, new_n_n904_,
    new_nw53_, new_n_n833_, new_n_n823_, new_n_n813_, new_nl55_, new_nv56_,
    new_n_n811_, new_n_n800_, new_n_n789_, new_n_n759_, new_n_n748_,
    new_n_n723_, new_n_n712_, new_n_n701_, new_n_n690_, new_n_n660_,
    new_n_n650_, new_n_n639_, new_n_n625_, new_n_n614_, new_n_n603_,
    new_n_n592_, new_n_n562_, new_n_n551_, new_n_n540_, new_n_n529_,
    new_n_n526_, new_n_n515_, new_n_n504_, new_n_n493_, new_n_n463_,
    new_n_n452_, new_n_n441_, new_n_n430_, new_n_n427_, new_n_n416_,
    new_n_n405_, new_n_n394_, new_n_n364_, new_n_n353_, new_n_n342_,
    new_n_n331_, new_n_n328_, new_n_n317_, new_n_n306_, new_n_n295_,
    new_n_n279_, new_n_n265_, new_n_n254_, new_n_n243_, new_n_n232_,
    new_n_n218_, new_n_n207_, new_n_n196_, new_n_n180_, new_n_n170_,
    new_n_n167_, new_n_n156_, new_n_n145_, new_n_n134_, new_n_n109_,
    new_n_n98_, new_nt5_, new_ni6_, new_nz6_, new_ni7_, new_nd8_,
    new_nl10_, new_nw10_, new_nq30_, new_n_n1147_, new_nu32_, new_nl33_,
    new_nu33_, new_nh34_, new_nq34_, new_nu35_, new_nd36_, new_nq36_,
    new_n_n1093_, new_n_n1090_, new_nk37_, new_ny37_, new_nl38_,
    new_n_n1063_, new_ne39_, new_nk39_, new_n_n1049_, new_ng40_, new_nl40_,
    new_nw40_, new_n_n1029_, new_nu41_, new_ny41_, new_n_n1011_, new_nm42_,
    new_nq42_, new_n_n994_, new_n_n962_, new_n_n958_, new_ni45_, new_nc47_,
    new_ni47_, new_nx53_, new_nf54_, new_n_n822_, new_n_n814_, new_nv55_,
    new_nw56_, new_nf57_, new_n_n799_, new_n_n790_, new_n_n758_,
    new_n_n749_, new_n_n722_, new_n_n713_, new_n_n700_, new_n_n691_,
    new_n_n659_, new_n_n651_, new_n_n629_, new_n_n624_, new_n_n615_,
    new_n_n602_, new_n_n593_, new_n_n561_, new_n_n552_, new_n_n539_,
    new_n_n530_, new_n_n525_, new_n_n516_, new_n_n503_, new_n_n494_,
    new_n_n462_, new_n_n453_, new_n_n440_, new_n_n431_, new_n_n426_,
    new_n_n417_, new_n_n404_, new_n_n395_, new_n_n363_, new_n_n354_,
    new_n_n341_, new_n_n332_, new_n_n327_, new_n_n318_, new_n_n305_,
    new_n_n296_, new_n_n269_, new_n_n264_, new_n_n255_, new_n_n242_,
    new_n_n233_, new_n_n228_, new_n_n206_, new_n_n197_, new_n_n179_,
    new_n_n171_, new_n_n166_, new_n_n157_, new_n_n144_, new_n_n135_,
    new_n_n108_, new_n_n99_, new_nu5_, new_nn6_, new_nw6_, new_nh7_,
    new_n_n1388_, new_nz9_, new_nc31_, new_nh31_, new_n_n1110_, new_nm33_,
    new_nx33_, new_ne34_, new_np34_, new_nv35_, new_ng36_, new_np36_,
    new_nb37_, new_ng37_, new_nl37_, new_n_n1079_, new_nk38_, new_n_n1070_,
    new_nz38_, new_ng39_, new_n_n1055_, new_ns39_, new_nf40_, new_n_n1046_,
    new_nq40_, new_ne41_, new_nt41_, new_n_n1015_, new_n_n1010_,
    new_n_n1007_, new_n_n1002_, new_nu42_, new_n_n964_, new_nj44_,
    new_n_n949_, new_ny53_, new_n_n831_, new_n_n825_, new_n_n815_,
    new_nf56_, new_nx56_, new_n_n809_, new_n_n802_, new_n_n791_,
    new_n_n739_, new_n_n728_, new_n_n721_, new_n_n710_, new_n_n703_,
    new_n_n692_, new_n_n658_, new_n_n641_, new_n_n630_, new_n_n623_,
    new_n_n612_, new_n_n605_, new_n_n594_, new_n_n560_, new_n_n549_,
    new_n_n542_, new_n_n531_, new_n_n524_, new_n_n513_, new_n_n506_,
    new_n_n495_, new_n_n479_, new_n_n461_, new_n_n450_, new_n_n443_,
    new_n_n432_, new_n_n425_, new_n_n414_, new_n_n407_, new_n_n396_,
    new_n_n380_, new_n_n369_, new_n_n362_, new_n_n351_, new_n_n344_,
    new_n_n333_, new_n_n326_, new_n_n315_, new_n_n308_, new_n_n297_,
    new_n_n281_, new_n_n270_, new_n_n263_, new_n_n252_, new_n_n245_,
    new_n_n234_, new_n_n227_, new_n_n216_, new_n_n198_, new_n_n182_,
    new_n_n172_, new_n_n165_, new_n_n154_, new_n_n147_, new_n_n136_,
    new_n_n129_, new_n_n118_, new_nv5_, new_nk6_, new_nx6_, new_ng7_,
    new_np7_, new_ny9_, new_n_n1140_, new_n_n1134_, new_n_n1104_,
    new_nn33_, new_nw33_, new_nf34_, new_no34_, new_nw35_, new_nf36_,
    new_n_n1098_, new_na37_, new_n_n1089_, new_n_n1083_, new_nq37_,
    new_nj38_, new_n_n1069_, new_nv38_, new_n_n1061_, new_n_n1056_,
    new_n_n1051_, new_ne40_, new_n_n1045_, new_n_n1039_, new_n_n1035_,
    new_n_n1022_, new_n_n1016_, new_na42_, new_nn42_, new_n_n1001_,
    new_n_n995_, new_n_n963_, new_n_n959_, new_ns44_, new_n_n839_,
    new_n_n832_, new_n_n824_, new_n_n816_, new_np56_, new_ny56_,
    new_n_n810_, new_n_n801_, new_n_n792_, new_n_n738_, new_n_n729_,
    new_n_n720_, new_n_n711_, new_n_n702_, new_n_n693_, new_n_n649_,
    new_n_n640_, new_n_n631_, new_n_n622_, new_n_n613_, new_n_n604_,
    new_n_n595_, new_n_n559_, new_n_n550_, new_n_n541_, new_n_n532_,
    new_n_n523_, new_n_n514_, new_n_n505_, new_n_n496_, new_n_n469_,
    new_n_n460_, new_n_n451_, new_n_n442_, new_n_n433_, new_n_n424_,
    new_n_n415_, new_n_n406_, new_n_n397_, new_n_n379_, new_n_n370_,
    new_n_n361_, new_n_n352_, new_n_n343_, new_n_n334_, new_n_n325_,
    new_n_n316_, new_n_n307_, new_n_n298_, new_n_n280_, new_n_n271_,
    new_n_n262_, new_n_n253_, new_n_n244_, new_n_n235_, new_n_n226_,
    new_n_n217_, new_n_n208_, new_n_n181_, new_n_n173_, new_n_n164_,
    new_n_n155_, new_n_n146_, new_n_n137_, new_n_n128_, new_n_n119_,
    new_nw5_, new_ni20_, new_n_n1347_, new_na21_, new_n_n1302_,
    new_n_n1293_, new_nv23_, new_n_n1280_, new_nj24_, new_n_n1269_,
    new_no25_, new_n_n1236_, new_n_n1229_, new_nk26_, new_n_n1219_,
    new_n_n1211_, new_n_n1206_, new_n_n1198_, new_nc28_, new_n_n1174_,
    new_n_n1167_, new_nr29_, new_nw29_, new_nc30_, new_nw30_, new_n_n1142_,
    new_n_n1135_, new_n_n1109_, new_n_n1103_, new_nr33_, new_nc34_,
    new_nn34_, new_np37_, new_ni38_, new_n_n84_, new_n_n73_, new_n_n62_,
    new_n_n51_, new_n_n40_, new_nk20_, new_n_n1348_, new_nn21_,
    new_n_n1301_, new_n_n1294_, new_n_n1287_, new_n_n1281_, new_nl24_,
    new_nq24_, new_n_n1243_, new_n_n1237_, new_n_n1228_, new_n_n1224_,
    new_n_n1218_, new_n_n1212_, new_n_n1205_, new_n_n1199_, new_ng28_,
    new_n_n1173_, new_n_n1168_, new_n_n1161_, new_n_n1155_, new_nd30_,
    new_nv30_, new_n_n1141_, new_ng31_, new_n_n1116_, new_n_n1102_,
    new_nq33_, new_nd34_, new_nm34_, new_n_n1080_, new_nh38_, new_n_n85_,
    new_n_n72_, new_n_n63_, new_n_n50_, new_n_n41_, new_ng20_, new_nq20_,
    new_n_n1331_, new_ne23_, new_ni23_, new_n_n1286_, new_n_n1279_,
    new_ng24_, new_n_n1270_, new_ns25_, new_ny25_, new_n_n1222_, new_nt26_,
    new_nz26_, new_no27_, new_nx27_, new_n_n1185_, new_n_n1172_,
    new_n_n1166_, new_nq29_, new_n_n1156_, new_nf30_, new_n_n1148_,
    new_nb31_, new_n_n1136_, new_n_n1117_, new_ng33_, new_nt33_, new_na34_,
    new_nl34_, new_n_n1092_, new_n_n1085_, new_n_n86_, new_n_n71_,
    new_n_n60_, new_n_n53_, new_n_n42_, new_nh20_, new_n_n1349_, new_na22_,
    new_n_n1303_, new_n_n1295_, new_nw23_, new_na24_, new_ni24_,
    new_n_n1271_, new_n_n1244_, new_n_n1227_, new_n_n1223_, new_nu26_,
    new_n_n1213_, new_n_n1197_, new_na28_, new_n_n1186_, new_nz28_,
    new_nf29_, new_n_n1162_, new_n_n1157_, new_nk30_, new_nx30_,
    new_n_n1143_, new_n_n1137_, new_n_n1123_, new_ni33_, new_ns33_,
    new_nb34_, new_nk34_, new_nf37_, new_n_n1086_, new_n_n87_, new_n_n70_,
    new_n_n61_, new_n_n52_, new_n_n43_, new_ns5_, new_nf10_, new_nt10_,
    new_nm16_, new_ne20_, new_n_n1350_, new_nm22_, new_n_n1305_,
    new_n_n1296_, new_nu24_, new_nx24_, new_n_n1249_, new_n_n1245_,
    new_n_n1226_, new_n_n1221_, new_n_n1216_, new_nj27_, new_n_n1201_,
    new_n_n1193_, new_nf28_, new_n_n1171_, new_n_n1165_, new_n_n1159_,
    new_nz29_, new_na30_, new_ns30_, new_n_n1144_, new_n_n1138_,
    new_n_n1122_, new_nh32_, new_nv32_, new_na33_, new_nj34_, new_ni36_,
    new_nr36_, new_nn47_, new_nw47_, new_n_n830_, new_n_n820_, new_n_n797_,
    new_n_n88_, new_n_n33_, new_n_n22_, new_n_n11_, new_n_n0_, new_nt6_,
    new_ne10_, new_nu10_, new_nj16_, new_nf20_, new_n_n1351_, new_n_n1323_,
    new_n_n1304_, new_ng23_, new_n_n1264_, new_n_n1257_, new_nc25_,
    new_nn25_, new_n_n1225_, new_nm26_, new_n_n1209_, new_nm27_, new_nq27_,
    new_n_n1192_, new_n_n1187_, new_n_n1170_, new_ng29_, new_n_n1158_,
    new_nx29_, new_nb30_, new_nr30_, new_nz30_, new_nf31_, new_nz31_,
    new_nf32_, new_n_n1113_, new_n_n1107_, new_nz33_, new_n_n1101_,
    new_n_n1096_, new_no47_, new_n_n900_, new_n_n829_, new_n_n821_,
    new_n_n807_, new_n_n89_, new_n_n32_, new_n_n23_, new_n_n10_, new_n_n1_,
    new_ne7_, new_nj10_, new_nr10_, new_n_n1380_, new_n_n1355_,
    new_n_n1352_, new_n_n1315_, new_n_n1263_, new_n_n1256_, new_n_n1251_,
    new_n_n1246_, new_na26_, new_nv26_, new_nd27_, new_n_n1207_, new_nr27_,
    new_nu27_, new_n_n1188_, new_nc29_, new_nh29_, new_n_n1160_,
    new_n_n1153_, new_n_n1150_, new_nu30_, new_ny30_, new_nd31_, new_nb32_,
    new_np32_, new_n_n1115_, new_n_n1108_, new_np33_, new_nn35_, new_ny35_,
    new_ng44_, new_nj47_, new_n_n901_, new_np53_, new_n_n837_, new_na57_,
    new_n_n31_, new_n_n20_, new_n_n13_, new_n_n2_, new_no7_, new_ng10_,
    new_ns10_, new_n_n1381_, new_nc20_, new_nn20_, new_n_n1306_,
    new_n_n1262_, new_nz24_, new_n_n1250_, new_n_n1247_, new_n_n1220_,
    new_n_n1217_, new_n_n1210_, new_nn27_, new_n_n1200_, new_n_n1194_,
    new_n_n1189_, new_n_n1169_, new_n_n1164_, new_ns29_, new_n_n1154_,
    new_n_n1149_, new_nt30_, new_n_n1145_, new_n_n1139_, new_nd32_,
    new_nl32_, new_n_n1114_, new_nz32_, new_nf33_, new_no35_, new_nx35_,
    new_nr44_, new_nl47_, new_nt47_, new_nq53_, new_n_n838_, new_nq56_,
    new_n_n30_, new_n_n21_, new_n_n12_, new_n_n3_, new_n_n1389_, new_nu16_,
    new_ne17_, new_nr17_, new_nc18_, new_n_n1344_, new_nd21_, new_n_n1334_,
    new_n_n1327_, new_ni22_, new_nu22_, new_n_n1317_, new_n_n1307_,
    new_n_n1278_, new_n_n1274_, new_n_n1267_, new_nw24_, new_n_n1252_,
    new_n_n1248_, new_n_n1238_, new_n_n1204_, new_n_n1196_, new_nd28_,
    new_nj28_, new_n_n1176_, new_no31_, new_nv31_, new_nt34_, new_ne35_,
    new_nz44_, new_nf48_, new_n_n892_, new_n_n886_, new_nr49_, new_nw52_,
    new_nc53_, new_ng56_, new_n_n59_, new_n_n48_, new_n_n37_, new_n_n26_,
    new_n_n15_, new_n_n4_, new_nc8_, new_n_n1378_, new_nd17_, new_n_n1368_,
    new_nb18_, new_n_n1343_, new_nc21_, new_n_n1333_, new_n_n1328_,
    new_nj22_, new_nt22_, new_n_n1316_, new_n_n1308_, new_nb24_, new_nm24_,
    new_n_n1266_, new_n_n1260_, new_nb25_, new_nm25_, new_n_n1232_,
    new_n_n1208_, new_n_n1195_, new_n_n1190_, new_n_n1179_, new_nu28_,
    new_n_n1132_, new_nt31_, new_nu34_, new_nd35_, new_ng45_, new_ng48_,
    new_n_n893_, new_nb49_, new_np49_, new_n_n847_, new_na53_, new_nw55_,
    new_n_n58_, new_n_n49_, new_n_n36_, new_n_n27_, new_n_n14_, new_n_n5_,
    new_nm8_, new_n_n1377_, new_ni17_, new_n_n1370_, new_n_n1363_,
    new_n_n1342_, new_nf21_, new_n_n1336_, new_n_n1329_, new_nk22_,
    new_n_n1324_, new_nc23_, new_n_n1309_, new_n_n1291_, new_n_n1284_,
    new_n_n1265_, new_n_n1258_, new_na25_, new_nl25_, new_n_n1240_,
    new_nw25_, new_nf27_, new_n_n1202_, new_n_n1191_, new_n_n1181_,
    new_nt28_, new_n_n1133_, new_n_n1127_, new_n_n938_, new_ni48_,
    new_n_n891_, new_nz48_, new_no49_, new_n_n856_, new_n_n853_, new_nm55_,
    new_n_n79_, new_n_n68_, new_n_n35_, new_n_n24_, new_n_n17_, new_n_n6_,
    new_nt8_, new_nw16_, new_nf17_, new_n_n1369_, new_n_n1364_,
    new_n_n1341_, new_ne21_, new_n_n1335_, new_n_n1330_, new_nl22_,
    new_nv22_, new_n_n1318_, new_n_n1310_, new_nt23_, new_n_n1285_,
    new_ns24_, new_n_n1259_, new_n_n1253_, new_nj25_, new_n_n1239_,
    new_nu25_, new_nh27_, new_n_n1203_, new_nt27_, new_n_n1180_, new_ns28_,
    new_nn31_, new_n_n1128_, new_n_n931_, new_nj48_, new_nq48_,
    new_n_n887_, new_nn49_, new_nc52_, new_n_n854_, new_nc55_, new_n_n78_,
    new_n_n69_, new_n_n34_, new_n_n25_, new_n_n16_, new_n_n7_, new_nd9_,
    new_nl18_, new_n_n1357_, new_nz19_, new_nr20_, new_n_n1338_, new_nr21_,
    new_nx21_, new_nc22_, new_nq22_, new_n_n1320_, new_n_n1311_,
    new_n_n1298_, new_nr23_, new_n_n1290_, new_nx23_, new_n_n1275_,
    new_n_n1272_, new_n_n1255_, new_ni25_, new_np25_, new_n_n1233_,
    new_nf26_, new_nr26_, new_n_n1214_, new_n_n1182_, new_nr28_, new_ns31_,
    new_n_n925_, new_nz49_, new_nl50_, new_n_n875_, new_np51_, new_n_n871_,
    new_n_n861_, new_ns54_, new_n_n80_, new_n_n77_, new_n_n66_, new_n_n55_,
    new_n_n44_, new_n_n19_, new_n_n8_, new_nn9_, new_nm18_, new_n_n1358_,
    new_nb20_, new_nt20_, new_n_n1339_, new_n_n1332_, new_nv21_, new_nd22_,
    new_np22_, new_n_n1319_, new_nd23_, new_n_n1297_, new_nq23_, new_nu23_,
    new_n_n1283_, new_nc24_, new_np24_, new_n_n1254_, new_ng25_, new_nr25_,
    new_n_n1234_, new_n_n1231_, new_ns26_, new_ny26_, new_ni28_, new_nq28_,
    new_nl31_, new_n_n918_, new_na50_, new_nj50_, new_n_n874_, new_nm51_,
    new_n_n870_, new_n_n862_, new_n_n812_, new_n_n81_, new_n_n76_,
    new_n_n67_, new_n_n54_, new_n_n45_, new_n_n18_, new_n_n9_, new_nx9_,
    new_np18_, new_ng19_, new_nv19_, new_n_n1354_, new_nv20_, new_nm21_,
    new_np21_, new_n_n1325_, new_nf22_, new_ns22_, new_nz22_, new_n_n1312_,
    new_n_n1300_, new_no23_, new_n_n1289_, new_n_n1282_, new_n_n1277_,
    new_n_n1273_, new_n_n1268_, new_n_n1261_, new_n_n1242_, new_n_n1235_,
    new_n_n1230_, new_nj26_, new_n_n1215_, new_n_n1184_, new_np28_,
    new_nr46_, new_n_n881_, new_np50_, new_nb51_, new_n_n872_, new_n_n82_,
    new_n_n75_, new_n_n64_, new_n_n57_, new_n_n46_, new_n_n39_, new_n_n28_,
    new_nq18_, new_ne19_, new_ny19_, new_n_n1346_, new_n_n1340_,
    new_n_n1337_, new_nq21_, new_n_n1326_, new_nh22_, new_nr22_,
    new_n_n1321_, new_n_n1313_, new_n_n1299_, new_n_n1292_, new_n_n1288_,
    new_nz23_, new_n_n1276_, new_no24_, new_nr24_, new_nv24_, new_n_n1241_,
    new_nt25_, new_nx25_, new_nh26_, new_no26_, new_n_n1183_, new_no28_,
    new_n_n908_, new_n_n880_, new_nn50_, new_nd51_, new_n_n873_,
    new_n_n83_, new_n_n74_, new_n_n65_, new_n_n56_, new_n_n47_, new_n_n38_,
    new_n_n29_;
  assign new_na1_ = pa1;
  assign new_nb2_ = pb2;
  assign new_nc3_ = pc3;
  assign new_nd4_ = pd4;
  assign new_ne5_ = pe5;
  assign pf6 = new_nf6_;
  assign pg7 = new_ng7_;
  assign ph8 = new_nh8_;
  assign pi9 = new_ni9_;
  assign new_np_ = pp;
  assign pq10 = new_nq10_;
  assign new_na0_ = pa0;
  assign new_nb3_ = pb3;
  assign new_nc2_ = pc2;
  assign new_nd5_ = pd5;
  assign new_ne4_ = pe4;
  assign pf7 = new_nf7_;
  assign pg6 = new_ng6_;
  assign ph9 = new_nh9_;
  assign pi8 = new_ni8_;
  assign pp10 = new_ng5_;
  assign new_nq_ = pq;
  assign new_na3_ = pa3;
  assign new_nb0_ = pb0;
  assign new_nc1_ = pc1;
  assign pd6 = new_nd6_;
  assign pe7 = new_ne7_;
  assign new_nf4_ = pf4;
  assign new_ng5_ = pg5;
  assign pj8 = new_nj8_;
  assign pk9 = new_nk9_;
  assign new_nr_ = pr;
  assign ps10 = new_ns10_;
  assign new_na2_ = pa2;
  assign new_nb1_ = pb1;
  assign new_nc0_ = pc0;
  assign pd7 = new_nd7_;
  assign pe6 = new_ne6_;
  assign new_nf5_ = pf5;
  assign new_ng4_ = pg4;
  assign pj9 = new_nj9_;
  assign pk8 = new_nk8_;
  assign pr10 = new_nr10_;
  assign new_ns_ = ps;
  assign new_na5_ = pa5;
  assign pb6 = new_nb6_;
  assign pc7 = new_nc7_;
  assign new_nd0_ = pd0;
  assign new_ne1_ = pe1;
  assign new_nf2_ = pf2;
  assign new_ng3_ = pg3;
  assign pl8 = new_nl8_;
  assign pm9 = new_nm9_;
  assign new_nt_ = pt;
  assign pu10 = new_nu10_;
  assign new_na4_ = pa4;
  assign pb7 = new_nb7_;
  assign pc6 = new_nc6_;
  assign new_nd1_ = pd1;
  assign new_ne0_ = pe0;
  assign new_nf3_ = pf3;
  assign new_ng2_ = pg2;
  assign pl9 = new_nl9_;
  assign pm8 = new_nm8_;
  assign pt10 = new_nt10_;
  assign new_nu_ = pu;
  assign pa7 = new_na7_;
  assign new_nb4_ = pb4;
  assign new_nc5_ = pc5;
  assign new_nd2_ = pd2;
  assign new_ne3_ = pe3;
  assign new_nf0_ = pf0;
  assign new_ng1_ = pg1;
  assign pn8 = new_nn8_;
  assign po9 = new_no9_;
  assign new_nv_ = pv;
  assign pw10 = new_nw10_;
  assign pa6 = new_na6_;
  assign new_nb5_ = pb5;
  assign new_nc4_ = pc4;
  assign new_nd3_ = pd3;
  assign new_ne2_ = pe2;
  assign new_nf1_ = pf1;
  assign new_ng0_ = pg0;
  assign pn9 = new_nn9_;
  assign po8 = new_no8_;
  assign pv10 = new_nv10_;
  assign new_nw_ = pw;
  assign pa9 = new_na9_;
  assign new_nh0_ = ph0;
  assign new_ni1_ = pi1;
  assign new_nj2_ = pj2;
  assign new_nk3_ = pk3;
  assign new_nl4_ = pl4;
  assign new_nm5_ = pm5;
  assign pn6 = new_nn6_;
  assign po7 = new_no7_;
  assign py10 = new_ny10_;
  assign pa8 = new_na8_;
  assign new_nh1_ = ph1;
  assign new_ni0_ = pi0;
  assign new_nj3_ = pj3;
  assign new_nk2_ = pk2;
  assign new_nl5_ = pl5;
  assign new_nm4_ = pm4;
  assign pn7 = new_nn7_;
  assign po6 = new_no6_;
  assign px10 = new_nx10_;
  assign new_ny_ = py;
  assign pb8 = new_nb8_;
  assign pc9 = new_nc9_;
  assign new_nh2_ = ph2;
  assign new_ni3_ = pi3;
  assign new_nj0_ = pj0;
  assign new_nk1_ = pk1;
  assign pl6 = new_na_;
  assign pm7 = new_nm7_;
  assign new_nn4_ = pn4;
  assign new_no5_ = po5;
  assign new_nz_ = pz;
  assign pb9 = new_nb9_;
  assign pc8 = new_nc8_;
  assign new_nh3_ = ph3;
  assign new_ni2_ = pi2;
  assign new_nj1_ = pj1;
  assign new_nk0_ = pk0;
  assign pl7 = new_nl7_;
  assign pm6 = new_ne1_;
  assign new_nn5_ = pn5;
  assign new_no4_ = po4;
  assign pd8 = new_nd8_;
  assign pe9 = new_ne9_;
  assign new_nh4_ = ph4;
  assign new_ni5_ = pi5;
  assign pj6 = new_nj6_;
  assign pk7 = new_nk7_;
  assign new_nl0_ = pl0;
  assign new_nm1_ = pm1;
  assign new_nn2_ = pn2;
  assign new_no3_ = po3;
  assign pd9 = new_nd9_;
  assign pe8 = new_ne8_;
  assign new_nh5_ = ph5;
  assign new_ni4_ = pi4;
  assign pj7 = new_nj7_;
  assign pk6 = new_nk6_;
  assign new_nl1_ = pl1;
  assign new_nm0_ = pm0;
  assign new_nn3_ = pn3;
  assign new_no2_ = po2;
  assign pf8 = new_nf8_;
  assign pg9 = new_ng9_;
  assign ph6 = new_nh6_;
  assign pi7 = new_ni7_;
  assign new_nj4_ = pj4;
  assign new_nk5_ = pk5;
  assign new_nl2_ = pl2;
  assign new_nm3_ = pm3;
  assign new_nn0_ = pn0;
  assign new_no1_ = po1;
  assign pf9 = new_nf9_;
  assign pg8 = new_ng8_;
  assign ph7 = new_nh7_;
  assign pi6 = new_ni6_;
  assign new_nj5_ = pj5;
  assign new_nk4_ = pk4;
  assign new_nl3_ = pl3;
  assign new_nm2_ = pm2;
  assign new_nn1_ = pn1;
  assign new_no0_ = po0;
  assign pa10 = new_na10_;
  assign new_np0_ = pp0;
  assign new_nq1_ = pq1;
  assign new_nr2_ = pr2;
  assign new_ns3_ = ps3;
  assign new_nt4_ = pt4;
  assign pu5 = new_nu5_;
  assign pv6 = new_nv6_;
  assign pw7 = new_nw7_;
  assign px8 = new_nx8_;
  assign py9 = new_ny9_;
  assign new_na_ = pa;
  assign new_np1_ = pp1;
  assign new_nq0_ = pq0;
  assign new_nr3_ = pr3;
  assign new_ns2_ = ps2;
  assign pt5 = new_nt5_;
  assign new_nu4_ = pu4;
  assign pv7 = new_nv7_;
  assign pw6 = new_nw6_;
  assign px9 = new_nx9_;
  assign py8 = new_ny8_;
  assign new_nb_ = pb;
  assign pc10 = new_nc10_;
  assign new_np2_ = pp2;
  assign new_nq3_ = pq3;
  assign new_nr0_ = pr0;
  assign new_ns1_ = ps1;
  assign pt6 = new_nt6_;
  assign pu7 = new_nu7_;
  assign new_nv4_ = pv4;
  assign pw5 = new_nw5_;
  assign pz8 = new_nz8_;
  assign pb10 = new_nb10_;
  assign new_nc_ = pc;
  assign new_np3_ = pp3;
  assign new_nq2_ = pq2;
  assign new_nr1_ = pr1;
  assign new_ns0_ = ps0;
  assign pt7 = new_nt7_;
  assign pu6 = new_nu6_;
  assign pv5 = new_nv5_;
  assign new_nw4_ = pw4;
  assign pz9 = new_nz9_;
  assign new_nd_ = pd;
  assign pe10 = new_ne10_;
  assign new_np4_ = pp4;
  assign new_nq5_ = pq5;
  assign pr6 = new_nj1_;
  assign ps7 = new_ns7_;
  assign new_nt0_ = pt0;
  assign new_nu1_ = pu1;
  assign new_nv2_ = pv2;
  assign new_nw3_ = pw3;
  assign pd10 = new_nd10_;
  assign new_ne_ = pe;
  assign new_np5_ = pp5;
  assign new_nq4_ = pq4;
  assign pr7 = new_nr7_;
  assign ps6 = new_ns6_;
  assign new_nt1_ = pt1;
  assign new_nu0_ = pu0;
  assign new_nv3_ = pv3;
  assign new_nw2_ = pw2;
  assign new_nf_ = pf;
  assign pg10 = new_ng10_;
  assign pp6 = new_np6_;
  assign pq7 = new_nq7_;
  assign new_nr4_ = pr4;
  assign ps5 = new_ns5_;
  assign new_nt2_ = pt2;
  assign new_nu3_ = pu3;
  assign new_nv0_ = pv0;
  assign new_nw1_ = pw1;
  assign pf10 = new_nf10_;
  assign new_ng_ = pg;
  assign pp7 = new_np7_;
  assign pq6 = new_nq6_;
  assign new_nr5_ = pr5;
  assign new_ns4_ = ps4;
  assign new_nt3_ = pt3;
  assign new_nu2_ = pu2;
  assign new_nv1_ = pv1;
  assign new_nw0_ = pw0;
  assign new_nh_ = ph;
  assign pi10 = new_na5_;
  assign pp8 = new_np8_;
  assign pq9 = new_nq9_;
  assign new_nx0_ = px0;
  assign new_ny1_ = py1;
  assign new_nz2_ = pz2;
  assign ph10 = new_ny_;
  assign new_ni_ = pi;
  assign pp9 = new_np9_;
  assign pq8 = new_nq8_;
  assign new_nx1_ = px1;
  assign new_ny0_ = py0;
  assign new_nz3_ = pz3;
  assign new_nj_ = pj;
  assign pk10 = new_nk10_;
  assign pr8 = new_nr8_;
  assign ps9 = new_ns9_;
  assign new_nx2_ = px2;
  assign new_ny3_ = py3;
  assign new_nz0_ = pz0;
  assign pj10 = new_nj10_;
  assign new_nk_ = pk;
  assign pr9 = new_nr9_;
  assign ps8 = new_ns8_;
  assign new_nx3_ = px3;
  assign new_ny2_ = py2;
  assign new_nz1_ = pz1;
  assign new_nl_ = pl;
  assign pm10 = new_nm10_;
  assign pt8 = new_nt8_;
  assign pu9 = new_nu9_;
  assign new_nx4_ = px4;
  assign py5 = new_ny5_;
  assign pz6 = new_nz6_;
  assign pl10 = new_nl10_;
  assign new_nm_ = pm;
  assign pt9 = new_nt9_;
  assign pu8 = new_nu8_;
  assign px5 = new_nx5_;
  assign new_ny4_ = py4;
  assign pz7 = new_nz7_;
  assign new_nn_ = pn;
  assign po10 = new_no10_;
  assign pv8 = new_nv8_;
  assign pw9 = new_nw9_;
  assign px6 = new_nx6_;
  assign py7 = new_ny7_;
  assign new_nz4_ = pz4;
  assign pn10 = new_nn10_;
  assign new_no_ = po;
  assign pv9 = new_nv9_;
  assign pw8 = new_nw8_;
  assign px7 = new_nx7_;
  assign py6 = new_ny6_;
  assign pz5 = new_nz5_;
  assign new_nf7_ = new_n_n268_ & new_n_n25_;
  assign new_nq7_ = new_nb_ | new_n_n35_;
  assign new_ny7_ = new_nt20_ & new_n_n47_;
  assign new_ng8_ = new_n_n57_ | new_n_n55_;
  assign new_n_n1384_ = new_n_n66_ & new_nj50_;
  assign new_nz8_ = new_n_n72_ | new_n_n76_;
  assign new_nk9_ = new_nz_ | new_n_n706_;
  assign new_nv9_ = new_nz_ | new_n_n97_;
  assign new_nj17_ = new_n_n136_ & new_n_n135_ & new_nu19_;
  assign new_nt17_ = new_n_n1365_ | new_n_n1366_;
  assign new_ne18_ = new_n_n1359_ | new_n_n1360_;
  assign new_nw18_ = new_n_n153_ | new_n_n152_;
  assign new_nq19_ = new_n_n159_ | new_n_n164_;
  assign new_n_n1314_ = new_n_n362_ & new_n_n201_ & new_nu22_;
  assign new_nb35_ = new_n_n398_ | new_n_n396_ | new_n_n397_ | new_n_n395_;
  assign new_nm35_ = new_n_n414_ | new_n_n447_;
  assign new_n_n1071_ = new_n_n520_ & new_n_n485_;
  assign new_n_n1064_ = new_n_n738_ & new_n_n490_;
  assign new_n_n1060_ = new_nj50_ & new_n_n492_;
  assign new_nn39_ = new_n_n1052_ | new_n_n1053_;
  assign new_n_n1047_ = new_n_n714_ & new_nw39_;
  assign new_n_n1024_ = new_nz50_ & new_nu3_;
  assign new_n_n1017_ = new_n_n533_ & new_n_n532_;
  assign new_ne42_ = new_n_n735_ & new_np41_;
  assign new_n_n1005_ = new_n_n563_ & new_n_n538_;
  assign new_n_n998_ = new_nz50_ & new_n_n542_;
  assign new_n_n991_ = new_n_n548_ & new_n_n547_;
  assign new_ne43_ = new_n_n736_ & new_nk42_;
  assign new_nm43_ = new_n_n978_ | new_n_n977_ | new_n_n976_;
  assign new_ni44_ = new_n_n959_ | new_n_n570_;
  assign new_nt44_ = new_n_n574_ | new_n_n573_;
  assign new_na45_ = new_n_n947_ | new_n_n946_ | new_n_n945_;
  assign new_n_n942_ = new_nl4_ & new_nk4_ & new_ng45_;
  assign new_ns45_ = new_n_n934_ | new_n_n933_ | new_n_n932_;
  assign new_ny45_ = new_nn4_ & new_nm4_ & new_nn45_;
  assign new_n_n920_ = new_n_n733_ & new_nb46_;
  assign new_n_n912_ = new_n_n594_ & new_n_n590_;
  assign new_n_n909_ = new_n_n595_ & new_n_n794_;
  assign new_n_n890_ = new_n_n609_ & new_n_n755_;
  assign new_n_n884_ = new_n_n611_ & new_n_n624_;
  assign new_nv49_ = new_n_n882_ | new_n_n883_;
  assign new_n_n877_ = new_n_n628_ & new_nx49_ & new_nf50_;
  assign new_nz50_ = new_n_n651_ & new_n_n635_;
  assign new_nl51_ = new_n_n872_ | new_n_n873_;
  assign new_nq51_ = new_n_n863_ | new_n_n862_ | new_n_n861_ | new_n_n860_ | new_n_n867_ | new_n_n865_ | new_n_n864_ | new_n_n866_ | new_n_n641_;
  assign new_n_n859_ = new_nm53_ & new_n_n645_;
  assign new_nj52_ = new_n_n710_ | new_nm53_ | new_n_n704_;
  assign new_n_n849_ = new_n_n672_ & new_nh40_;
  assign new_n_n841_ = new_n_n657_ & new_n_n709_ & new_n_n672_;
  assign new_no53_ = new_nh40_ | new_no49_ | new_n_n687_;
  assign new_nl54_ = new_n_n683_ | new_n_n781_;
  assign new_nw54_ = new_n_n696_ | new_n_n694_ | new_n_n695_ | new_n_n693_;
  assign new_nh55_ = new_n_n712_ | new_n_n795_;
  assign new_ns55_ = new_n_n733_ | new_n_n787_;
  assign new_nd56_ = new_n_n754_ | new_n_n779_;
  assign new_no56_ = new_n_n765_ | new_n_n766_ | new_n_n767_;
  assign new_nz56_ = new_n_n794_ | new_n_n793_;
  assign new_n_n785_ = ~new_nr0_;
  assign new_n_n774_ = ~new_nj56_;
  assign new_n_n763_ = ~new_no3_;
  assign new_n_n752_ = ~new_nq56_;
  assign new_n_n741_ = ~new_nx55_;
  assign new_n_n730_ = ~new_nx4_;
  assign new_n_n719_ = ~new_na55_;
  assign new_n_n708_ = ~new_nm4_;
  assign new_n_n686_ = ~new_nq5_;
  assign new_n_n675_ = ~new_nb0_;
  assign new_n_n664_ = ~new_nh53_;
  assign new_n_n654_ = ~new_nq51_;
  assign new_n_n643_ = ~new_np50_;
  assign new_n_n632_ = ~new_ne0_;
  assign new_n_n621_ = ~new_na51_;
  assign new_n_n610_ = ~new_ny47_;
  assign new_n_n599_ = ~new_ni47_;
  assign new_n_n588_ = ~new_ng46_;
  assign new_n_n577_ = ~new_ni44_;
  assign new_n_n566_ = ~new_nv43_;
  assign new_n_n555_ = ~new_nl43_;
  assign new_n_n544_ = ~new_nv42_;
  assign new_n_n533_ = ~new_no41_;
  assign new_n_n522_ = ~new_nz40_;
  assign new_n_n511_ = ~new_ne39_;
  assign new_n_n500_ = ~new_nn39_;
  assign new_n_n489_ = ~new_ni38_;
  assign new_n_n478_ = ~new_no37_;
  assign new_n_n467_ = ~new_nz36_;
  assign new_n_n456_ = ~new_nt35_;
  assign new_n_n445_ = ~new_np_;
  assign new_n_n434_ = ~new_nd1_;
  assign new_n_n423_ = ~new_nh35_;
  assign new_n_n412_ = ~new_nw1_;
  assign new_n_n401_ = ~new_nv34_;
  assign new_n_n390_ = ~new_ny2_;
  assign new_n_n368_ = ~new_nj34_;
  assign new_n_n357_ = ~new_na1_;
  assign new_n_n346_ = ~new_nm33_;
  assign new_n_n335_ = ~new_nz0_;
  assign new_n_n324_ = ~new_ne19_;
  assign new_n_n313_ = ~new_ne32_;
  assign new_n_n302_ = ~new_nv31_;
  assign new_n_n291_ = ~new_nx30_;
  assign new_n_n258_ = ~new_nj27_;
  assign new_n_n247_ = ~new_nl_;
  assign new_n_n236_ = ~new_nr25_;
  assign new_n_n225_ = ~new_na25_;
  assign new_n_n214_ = ~new_ns24_;
  assign new_n_n203_ = ~new_ng23_;
  assign new_n_n192_ = ~new_nl22_;
  assign new_n_n149_ = ~new_ng1_;
  assign new_n_n138_ = ~new_ni17_;
  assign new_n_n127_ = ~new_nu19_;
  assign new_n_n116_ = ~new_na50_;
  assign new_n_n105_ = ~new_nt47_;
  assign new_n_n94_ = ~new_nv45_;
  assign new_nu6_ = new_n_n268_ & new_nx21_;
  assign new_nr7_ = new_nb_ | new_n_n36_;
  assign new_nx7_ = new_nt20_ & new_n_n46_;
  assign new_nh8_ = new_n_n57_ | new_n_n56_;
  assign new_nq8_ = new_n_n1384_ | new_n_n1383_ | new_n_n1382_;
  assign new_na9_ = new_n_n72_ | new_n_n77_;
  assign new_nj9_ = new_nz_ | new_n_n86_;
  assign new_nw9_ = new_n_n101_ & new_n_n99_ & new_n_n98_ & new_n_n100_;
  assign new_nl17_ = new_n_n136_ & new_na1_ & new_nu19_ & new_nz0_;
  assign new_n_n1367_ = new_n_n139_ & new_n_n382_;
  assign new_n_n1360_ = new_n_n142_ & new_nu18_;
  assign new_nu18_ = new_n_n151_ | new_n_n163_;
  assign new_nu19_ = new_nj18_ | new_n_n160_;
  assign new_n_n1322_ = new_n_n362_ & new_n_n338_;
  assign new_nc35_ = new_n_n402_ | new_n_n400_ | new_n_n401_ | new_n_n399_;
  assign new_nl35_ = new_n_n413_ | new_n_n445_;
  assign new_nq38_ = new_n_n1069_ | new_n_n1070_;
  assign new_n_n1065_ = new_nn3_ & new_nv38_;
  assign new_n_n1059_ = new_n_n520_ & new_n_n493_;
  assign new_n_n1054_ = new_n_n520_ & new_n_n498_;
  assign new_nk40_ = new_nt3_ & new_nr3_ & new_n_n511_ & new_ns3_;
  assign new_n_n1023_ = new_n_n563_ & new_n_n734_;
  assign new_nx41_ = new_n_n1017_ | new_n_n1016_ | new_n_n1015_;
  assign new_ng42_ = new_nr41_ & new_nx3_;
  assign new_n_n1006_ = new_nz50_ & new_n_n537_;
  assign new_n_n997_ = new_n_n563_ & new_n_n543_;
  assign new_nx42_ = new_n_n991_ | new_n_n990_ | new_n_n989_;
  assign new_ng43_ = new_nm42_ & new_na4_;
  assign new_n_n979_ = new_n_n736_ & new_nn43_;
  assign new_nv43_ = new_n_n963_ | new_n_n964_;
  assign new_nv44_ = new_n_n953_ | new_n_n954_;
  assign new_n_n948_ = new_n_n707_ & new_n_n578_;
  assign new_no45_ = new_n_n940_ | new_n_n941_;
  assign new_n_n935_ = new_n_n757_ & new_ng45_;
  assign new_nb46_ = new_nn45_ & new_nm4_;
  assign new_n_n921_ = new_nn4_ & new_n_n587_;
  assign new_np46_ = new_n_n591_ | new_n_n684_ | new_n_n592_;
  assign new_nx46_ = new_n_n909_ | new_n_n908_ | new_n_n907_;
  assign new_ns48_ = new_n_n782_ | new_ny47_;
  assign new_n_n885_ = new_n_n611_ & new_nr49_;
  assign new_n_n883_ = new_nr49_ & new_n_n657_;
  assign new_n_n878_ = new_n_n630_ & new_n_n628_ & new_nf50_;
  assign new_na51_ = new_ni5_ | new_n_n636_;
  assign new_nk51_ = new_n_n704_ & new_nl50_;
  assign new_n_n867_ = new_n_n686_ & new_n_n711_ & new_n_n710_;
  assign new_nv51_ = new_n_n858_ | new_n_n859_;
  assign new_nk52_ = new_n_n654_ & new_nv10_;
  assign new_n_n850_ = new_n_n672_ & new_no49_;
  assign new_n_n840_ = new_nh40_ & new_n_n709_ & new_n_n672_;
  assign new_nn53_ = new_no49_ | new_n_n669_;
  assign new_nm54_ = new_nc52_ | new_n_n783_;
  assign new_nv54_ = new_n_n690_ | new_n_n691_ | new_n_n692_;
  assign new_ni55_ = new_n_n713_ | new_n_n797_;
  assign new_nr55_ = new_n_n732_ | new_n_n785_;
  assign new_ne56_ = new_n_n755_ | new_n_n781_;
  assign new_nn56_ = new_n_n764_ | new_n_n799_;
  assign new_n_n808_ = ~new_nw56_;
  assign new_n_n784_ = ~new_ni4_;
  assign new_n_n775_ = ~new_nk56_;
  assign new_n_n762_ = ~new_nh3_;
  assign new_n_n753_ = ~new_np56_;
  assign new_n_n740_ = ~new_nw55_;
  assign new_n_n731_ = ~new_ne4_;
  assign new_n_n718_ = ~new_nz54_;
  assign new_n_n709_ = ~new_nm5_;
  assign new_n_n685_ = ~new_nn5_;
  assign new_n_n676_ = ~new_nz_;
  assign new_n_n663_ = ~new_ng53_;
  assign new_nv10_ = ~new_nu53_;
  assign new_n_n642_ = ~new_nr50_;
  assign new_n_n633_ = ~new_nt50_;
  assign new_n_n620_ = ~new_nt49_;
  assign new_n_n611_ = ~new_ny48_;
  assign new_n_n589_ = ~new_ny45_;
  assign new_n_n587_ = ~new_nb46_;
  assign new_n_n578_ = ~new_nn44_;
  assign new_n_n565_ = ~new_ny43_;
  assign new_n_n556_ = ~new_nk43_;
  assign new_n_n543_ = ~new_ng42_;
  assign new_n_n534_ = ~new_na42_;
  assign new_n_n521_ = ~new_nj40_;
  assign new_n_n512_ = ~new_nn40_;
  assign new_n_n499_ = ~new_nq39_;
  assign new_n_n490_ = ~new_nv38_;
  assign new_n_n488_ = ~new_nh38_;
  assign new_n_n466_ = ~new_nh0_;
  assign new_n_n457_ = ~new_nu35_;
  assign new_n_n444_ = ~new_nx1_;
  assign new_n_n435_ = ~new_nu_;
  assign new_n_n422_ = ~new_ng35_;
  assign new_n_n413_ = ~new_nz1_;
  assign new_n_n400_ = ~new_nu34_;
  assign new_n_n391_ = ~new_nc3_;
  assign new_n_n367_ = ~new_ni34_;
  assign new_n_n358_ = ~new_nb2_;
  assign new_n_n345_ = ~new_nl33_;
  assign new_n_n336_ = ~new_ne2_;
  assign new_n_n323_ = ~new_ny32_;
  assign new_n_n314_ = ~new_nd32_;
  assign new_n_n301_ = ~new_nv30_;
  assign new_n_n292_ = ~new_nr30_;
  assign new_n_n268_ = ~new_nb_;
  assign new_n_n246_ = ~new_nh26_;
  assign new_n_n237_ = ~new_nv19_;
  assign new_n_n224_ = ~new_nc25_;
  assign new_n_n215_ = ~new_nq24_;
  assign new_n_n202_ = ~new_nu22_;
  assign new_n_n193_ = ~new_nm22_;
  assign new_n_n148_ = ~new_ne1_;
  assign new_n_n139_ = ~new_nl17_;
  assign new_n_n126_ = ~new_nh54_;
  assign new_n_n117_ = ~new_nc50_;
  assign new_n_n104_ = ~new_nr47_;
  assign new_n_n95_ = ~new_ne46_;
  assign new_nf6_ = new_n_n8_ & new_n_n3_;
  assign new_nh6_ = new_n_n8_ & new_n_n5_;
  assign new_ns7_ = new_nb_ | new_n_n37_;
  assign new_na8_ = new_n_n57_ | new_n_n49_;
  assign new_ne8_ = new_nt20_ & new_n_n53_;
  assign new_np8_ = new_n_n72_ | new_n_n65_;
  assign new_nb9_ = new_n_n676_ & new_n_n78_;
  assign new_nm9_ = new_nz_ | new_n_n88_;
  assign new_nt9_ = new_nz_ | new_n_n95_;
  assign new_no16_ = new_nv0_ & new_nw0_ & new_nu19_;
  assign new_n_n1375_ = new_n_n131_ & new_n_n406_;
  assign new_n_n1359_ = new_n_n142_ & new_n_n155_;
  assign new_ny18_ = new_n_n1357_ | new_n_n1358_;
  assign new_nm19_ = new_n_n335_ & new_nk19_;
  assign new_nn22_ = new_nn1_ | new_n_n196_;
  assign new_n_n1129_ = new_n_n300_ & new_n_n301_;
  assign new_nz34_ = new_n_n391_ | new_n_n451_;
  assign new_nk35_ = new_n_n412_ | new_n_n443_;
  assign new_n_n1073_ = new_n_n485_ & new_n_n484_;
  assign new_nu38_ = new_n_n1064_ | new_n_n1065_;
  assign new_nh39_ = new_n_n1057_ | new_n_n1058_;
  assign new_nt39_ = new_n_n1047_ | new_n_n1048_;
  assign new_nj40_ = new_ns3_ & new_nr3_ & new_n_n510_;
  assign new_n_n1025_ = new_nw3_ & new_nv3_ & new_nu3_;
  assign new_nv41_ = new_n_n568_ & new_n_n531_;
  assign new_nh42_ = new_np41_ & new_n_n735_ & new_n_n760_;
  assign new_n_n1004_ = new_nx3_ & new_n_n539_;
  assign new_ns42_ = new_n_n999_ | new_n_n998_ | new_n_n997_;
  assign new_nv42_ = new_n_n568_ & new_n_n546_;
  assign new_nq43_ = new_n_n971_ | new_n_n972_;
  assign new_n_n965_ = new_n_n563_ & new_n_n564_;
  assign new_n_n954_ = new_ng4_ & new_n_n591_;
  assign new_n_n946_ = new_nv50_ & new_n_n759_;
  assign new_nk45_ = new_ng45_ & new_nk4_;
  assign new_n_n936_ = new_nk4_ & new_n_n581_;
  assign new_nd46_ = new_n_n925_ | new_n_n926_;
  assign new_n_n919_ = new_n_n588_ & new_n_n736_;
  assign new_n_n914_ = new_n_n590_ & new_n_n761_;
  assign new_n_n910_ = new_n_n788_ & new_nu46_;
  assign new_n_n899_ = new_nn47_ & new_nu4_;
  assign new_n_n896_ = new_n_n606_ & new_n_n683_;
  assign new_n_n882_ = new_n_n625_ & new_no49_;
  assign new_nf50_ = new_nt50_ & new_n_n656_;
  assign new_nv50_ = new_n_n633_ | new_n_n638_;
  assign new_nj51_ = new_nl5_ & new_n_n685_ & new_n_n676_ & new_n_n709_;
  assign new_n_n869_ = new_n_n704_ & new_nr5_ & new_nf52_;
  assign new_nu51_ = new_nj5_ & new_n_n646_;
  assign new_nl52_ = new_n_n682_ & new_n_n685_ & new_n_n676_ & new_nm5_;
  assign new_nv52_ = new_n_n682_ & new_nn5_ & new_n_n676_ & new_n_n709_;
  assign new_n_n843_ = new_nh40_ & new_n_n685_ & new_n_n672_;
  assign new_nm53_ = new_n_n668_ | new_n_n667_;
  assign new_nj54_ = new_n_n681_ & new_n_n680_ & new_n_n679_;
  assign new_nu54_ = new_n_n689_ | new_n_n799_;
  assign new_nj55_ = new_n_n714_ | new_n_n799_;
  assign new_nu55_ = new_n_n735_ | new_n_n791_;
  assign new_nb56_ = new_n_n750_ | new_n_n748_ | new_n_n749_ | new_n_n747_;
  assign new_nm56_ = new_n_n763_ | new_n_n797_;
  assign new_n_n798_ = ~new_np3_;
  assign new_n_n787_ = ~new_nq0_;
  assign new_n_n776_ = ~new_nd57_;
  assign new_n_n761_ = ~new_nb4_;
  assign new_n_n750_ = ~new_nv55_;
  assign new_n_n743_ = ~new_no55_;
  assign new_n_n732_ = ~new_nj4_;
  assign new_n_n699_ = ~new_nq54_;
  assign new_n_n688_ = ~new_nl3_;
  assign new_n_n677_ = ~new_nw53_;
  assign new_n_n662_ = ~new_nf53_;
  assign new_n_n652_ = ~new_ng49_;
  assign new_n_n645_ = ~new_nj5_;
  assign new_n_n634_ = ~new_nd47_;
  assign new_n_n619_ = ~new_nj10_;
  assign new_n_n601_ = ~new_nn47_;
  assign new_n_n590_ = ~new_nj46_;
  assign new_n_n564_ = ~new_nj43_;
  assign new_n_n553_ = ~new_nm42_;
  assign new_n_n546_ = ~new_ns42_;
  assign new_n_n535_ = ~new_ny41_;
  assign new_n_n520_ = ~new_nj50_;
  assign new_n_n509_ = ~new_nb39_;
  assign new_n_n502_ = ~new_nz38_;
  assign new_n_n491_ = ~new_nt38_;
  assign new_n_n465_ = ~new_no36_;
  assign new_n_n454_ = ~new_nc36_;
  assign new_n_n447_ = ~new_no_;
  assign new_n_n436_ = ~new_ng2_;
  assign new_n_n421_ = ~new_nf35_;
  assign new_n_n410_ = ~new_nm2_;
  assign new_n_n403_ = ~new_np35_;
  assign new_n_n392_ = ~new_nx34_;
  assign new_n_n366_ = ~new_nb3_;
  assign new_n_n355_ = ~new_nm34_;
  assign new_n_n348_ = ~new_no33_;
  assign new_n_n337_ = ~new_nn1_;
  assign new_n_n322_ = ~new_nz32_;
  assign new_n_n311_ = ~new_nl31_;
  assign new_n_n304_ = ~new_nr31_;
  assign new_n_n293_ = ~new_np30_;
  assign new_n_n267_ = ~new_nn2_;
  assign new_n_n256_ = ~new_nf27_;
  assign new_n_n238_ = ~new_nl25_;
  assign new_n_n223_ = ~new_nj24_;
  assign new_n_n212_ = ~new_nt23_;
  assign new_n_n205_ = ~new_nv23_;
  assign new_n_n194_ = ~new_ne21_;
  assign new_n_n169_ = ~new_ni19_;
  assign new_n_n158_ = ~new_ng_;
  assign new_n_n125_ = ~new_ng54_;
  assign new_n_n114_ = ~new_nm49_;
  assign new_n_n107_ = ~new_nj48_;
  assign new_n_n96_ = ~new_nh46_;
  assign new_ng6_ = new_n_n8_ & new_n_n4_;
  assign new_nt7_ = new_nb_ | new_n_n38_;
  assign new_nz7_ = new_nt20_ & new_n_n48_;
  assign new_nf8_ = new_nt20_ & new_n_n54_;
  assign new_no8_ = new_ne52_ & new_n_n64_;
  assign new_nc9_ = new_n_n676_ & new_n_n79_;
  assign new_nl9_ = new_nz_ | new_n_n87_;
  assign new_nu9_ = new_nz_ | new_n_n96_;
  assign new_nq16_ = new_nv0_ & new_nx0_ & new_nu19_ & new_nw0_;
  assign new_n_n1376_ = new_no16_ & new_nx0_;
  assign new_nj18_ = new_nh1_ | new_n_n143_;
  assign new_nx18_ = new_n_n154_ & new_n_n155_;
  assign new_no19_ = new_nb_ | new_nm1_ | new_n_n334_ | new_n_n337_;
  assign new_nb22_ = new_n_n341_ | new_nh22_;
  assign new_ny31_ = new_n_n1122_ | new_n_n1123_;
  assign new_na35_ = new_n_n392_ | new_n_n393_ | new_n_n394_;
  assign new_nj35_ = new_n_n411_ | new_n_n441_;
  assign new_n_n1072_ = new_nj50_ & new_n_n484_;
  assign new_n_n1066_ = new_n_n520_ & new_n_n489_;
  assign new_n_n1053_ = new_np3_ & new_n_n499_;
  assign new_n_n1048_ = new_nq3_ & new_n_n504_;
  assign new_ni40_ = new_n_n509_ & new_n_n739_ & new_n_n764_;
  assign new_ns41_ = new_n_n1023_ | new_n_n1024_;
  assign new_n_n1018_ = new_n_n567_ & new_n_n713_;
  assign new_nj42_ = new_ny3_ & new_nx3_ & new_nr41_;
  assign new_no42_ = new_n_n1003_ | new_n_n1004_;
  assign new_n_n999_ = new_n_n543_ & new_n_n542_;
  assign new_n_n992_ = new_n_n567_ & new_n_n798_;
  assign new_n_n972_ = new_nb4_ & new_n_n559_;
  assign new_n_n966_ = new_nz50_ & new_n_n562_;
  assign new_n_n953_ = new_n_n684_ & new_nt44_;
  assign new_n_n947_ = new_n_n576_ & new_n_n759_;
  assign new_nn45_ = new_n_n942_ | new_nj0_;
  assign new_nr45_ = new_n_n935_ | new_n_n936_;
  assign new_n_n926_ = new_nm4_ & new_n_n585_;
  assign new_nh46_ = new_n_n919_ | new_n_n918_ | new_n_n917_;
  assign new_n_n913_ = new_nv50_ & new_n_n761_;
  assign new_n_n911_ = new_nq4_ & new_n_n593_;
  assign new_n_n898_ = new_n_n601_ & new_n_n780_;
  assign new_n_n897_ = new_nj47_ & new_nv4_;
  assign new_nx49_ = new_nh5_ | new_n_n626_;
  assign new_n_n876_ = new_n_n630_ & new_n_n629_ & new_nf50_;
  assign new_ny50_ = new_ng49_ | new_n_n634_;
  assign new_ni51_ = new_n_n653_ & new_nv10_;
  assign new_n_n868_ = new_n_n704_ & new_nr5_ & new_nu53_;
  assign new_n_n860_ = new_n_n644_ & new_n_n643_ & new_n_n642_;
  assign new_nm52_ = new_n_n854_ | new_n_n853_ | new_n_n852_;
  assign new_n_n848_ = new_n_n672_ & new_n_n687_;
  assign new_n_n842_ = new_nm53_ & new_n_n709_ & new_n_n672_;
  assign new_nk53_ = new_n_n665_ | new_nj51_ | new_n_n666_;
  assign new_nk54_ = new_n_n682_ | new_n_n779_;
  assign new_nt54_ = new_n_n688_ | new_n_n797_;
  assign new_nk55_ = new_n_n715_ | new_n_n716_ | new_n_n717_;
  assign new_nt55_ = new_n_n734_ | new_n_n789_;
  assign new_nc56_ = new_n_n753_ & new_n_n752_ & new_n_n751_;
  assign new_nl56_ = new_n_n762_ | new_n_n795_;
  assign new_n_n788_ = ~new_nq4_;
  assign new_n_n786_ = ~new_nl4_;
  assign new_n_n777_ = ~new_nf57_;
  assign new_n_n760_ = ~new_ny3_;
  assign new_n_n751_ = ~new_no56_;
  assign new_n_n742_ = ~new_ny55_;
  assign new_n_n733_ = ~new_nn4_;
  assign new_n_n698_ = ~new_np54_;
  assign new_n_n689_ = ~new_nh40_;
  assign new_n_n687_ = ~new_nk40_;
  assign new_n_n661_ = ~new_nu52_;
  assign new_n_n653_ = ~new_np49_;
  assign new_n_n644_ = ~new_nn50_;
  assign new_n_n635_ = ~new_ng0_;
  assign new_n_n609_ = ~new_ng48_;
  assign new_n_n600_ = ~new_nl47_;
  assign new_n_n591_ = ~new_nt44_;
  assign new_n_n563_ = ~new_nz50_;
  assign new_n_n554_ = ~new_nn43_;
  assign new_n_n545_ = ~new_nt42_;
  assign new_n_n536_ = ~new_nx41_;
  assign new_n_n519_ = ~new_ni40_;
  assign new_n_n510_ = ~new_nd39_;
  assign new_n_n501_ = ~new_nm39_;
  assign new_n_n492_ = ~new_nj38_;
  assign new_n_n464_ = ~new_na37_;
  assign new_n_n455_ = ~new_nd36_;
  assign new_n_n446_ = ~new_na2_;
  assign new_n_n437_ = ~new_nt_;
  assign new_n_n420_ = ~new_ne35_;
  assign new_n_n411_ = ~new_nt1_;
  assign new_n_n402_ = ~new_nw34_;
  assign new_n_n393_ = ~new_ny34_;
  assign new_n_n365_ = ~new_nx2_;
  assign new_n_n356_ = ~new_nv0_;
  assign new_n_n347_ = ~new_nn33_;
  assign new_n_n338_ = ~new_nq1_;
  assign new_n_n321_ = ~new_nc33_;
  assign new_n_n312_ = ~new_nh32_;
  assign new_n_n303_ = ~new_ns31_;
  assign new_n_n294_ = ~new_nd31_;
  assign new_n_n266_ = ~new_nt26_;
  assign new_n_n257_ = ~new_nq27_;
  assign new_n_n248_ = ~new_nr26_;
  assign new_n_n222_ = ~new_nl24_;
  assign new_n_n213_ = ~new_nr23_;
  assign new_n_n204_ = ~new_nx23_;
  assign new_n_n195_ = ~new_nj22_;
  assign new_n_n168_ = ~new_nk19_;
  assign new_n_n159_ = ~new_no19_;
  assign new_n_n124_ = ~new_nf54_;
  assign new_n_n115_ = ~new_nn49_;
  assign new_n_n106_ = ~new_nw47_;
  assign new_n_n97_ = ~new_nk46_;
  assign new_nd6_ = new_n_n8_ & new_n_n1_;
  assign new_nu7_ = new_n_n42_ & new_n_n40_ & new_n_n39_ & new_n_n41_;
  assign new_n_n1387_ = new_n_n328_ & new_ne19_;
  assign new_nk8_ = new_n_n57_ | new_n_n60_;
  assign new_ns8_ = new_ne52_ & new_n_n68_;
  assign new_nv8_ = new_n_n72_ | new_n_n71_;
  assign new_ng9_ = new_nz_ | new_n_n83_;
  assign new_nr9_ = new_nz_ | new_n_n93_;
  assign new_nr16_ = new_n_n1379_ | new_nl16_;
  assign new_n_n1374_ = new_nq16_ & new_ny0_;
  assign new_n_n1371_ = new_n_n137_ & new_n_n335_;
  assign new_ny17_ = new_n_n1363_ | new_n_n1364_;
  assign new_ni19_ = new_nm19_ & new_n_n382_ & new_n_n407_ & new_n_n357_;
  assign new_nt21_ = new_n_n1329_ | new_n_n1327_ | new_n_n1326_ | new_n_n1325_ | new_n_n1328_ | new_n_n1330_;
  assign new_n_n1131_ = new_n_n301_ & new_ne19_;
  assign new_n_n1124_ = new_n_n305_ & new_n_n306_;
  assign new_nx34_ = new_n_n389_ | new_n_n447_;
  assign new_ni35_ = new_n_n410_ | new_n_n439_;
  assign new_nn38_ = new_nc52_ & new_n_n483_;
  assign new_n_n1067_ = new_nj50_ & new_n_n488_;
  assign new_nn40_ = new_nc52_ & new_n_n513_;
  assign new_nv40_ = new_n_n1036_ | new_n_n1035_ | new_n_n1034_;
  assign new_n_n1030_ = new_n_n734_ & new_n_n568_;
  assign new_nk42_ = new_n_n1009_ | new_ni0_;
  assign new_np42_ = new_n_n1002_ | new_n_n1001_ | new_n_n1000_;
  assign new_n_n986_ = new_n_n550_ & new_n_n714_;
  assign new_n_n981_ = new_n_n563_ & new_n_n553_;
  assign new_n_n974_ = new_nz50_ & new_n_n557_;
  assign new_n_n967_ = new_n_n564_ & new_n_n562_;
  assign new_nw44_ = new_n_n952_ | new_n_n951_ | new_n_n950_;
  assign new_ne45_ = new_n_n943_ | new_n_n944_;
  assign new_np45_ = new_n_n939_ | new_n_n938_ | new_n_n937_;
  assign new_nu45_ = new_n_n930_ | new_n_n931_;
  assign new_nv45_ = new_n_n929_ | new_n_n928_ | new_n_n927_;
  assign new_n_n923_ = new_nv50_ & new_n_n792_;
  assign new_n_n915_ = new_n_n758_ & new_ny45_;
  assign new_nw46_ = new_n_n910_ | new_n_n911_;
  assign new_ny47_ = new_n_n603_ | new_n_n602_;
  assign new_n_n895_ = new_nf48_ & new_nw4_;
  assign new_n_n888_ = new_n_n610_ & new_nz4_;
  assign new_nm49_ = new_no49_ | new_n_n614_ | new_n_n615_;
  assign new_nr50_ = new_n_n683_ & new_np50_;
  assign new_ng51_ = new_nl50_ & new_nr4_;
  assign new_n_n864_ = new_n_n686_ & new_n_n644_ & new_n_n643_;
  assign new_n_n857_ = new_nu51_ & new_nk5_;
  assign new_ne52_ = new_n_n669_ & new_n_n676_;
  assign new_nt52_ = new_nl5_ & new_nn5_ & new_n_n676_ & new_nm5_;
  assign new_n_n845_ = new_nm53_ & new_n_n685_ & new_n_n672_;
  assign new_ni53_ = new_n_n664_ & new_n_n669_ & new_n_n674_;
  assign new_np54_ = new_n_n685_ | new_n_n789_;
  assign new_na55_ = new_n_n705_ | new_n_n781_;
  assign new_nd55_ = new_n_n708_ | new_n_n787_;
  assign new_no55_ = new_n_n729_ | new_n_n779_;
  assign new_nz55_ = new_n_n740_ | new_n_n741_ | new_n_n742_;
  assign new_nk56_ = new_n_n761_ | new_n_n793_;
  assign new_n_n781_ = ~new_nt0_;
  assign new_n_n770_ = ~new_nf56_;
  assign new_n_n767_ = ~new_nn56_;
  assign new_n_n756_ = ~new_nf4_;
  assign new_n_n745_ = ~new_nq55_;
  assign new_n_n734_ = ~new_nu3_;
  assign new_n_n682_ = ~new_nl5_;
  assign new_n_n671_ = ~new_nv53_;
  assign new_n_n657_ = ~new_no49_;
  assign new_n_n647_ = ~new_nu51_;
  assign new_n_n636_ = ~new_no5_;
  assign new_n_n584_ = ~new_nu45_;
  assign new_n_n573_ = ~new_nr44_;
  assign new_n_n548_ = ~new_nj42_;
  assign new_n_n537_ = ~new_np41_;
  assign new_n_n485_ = ~new_nf38_;
  assign new_n_n474_ = ~new_np36_;
  assign new_n_n438_ = ~new_nj2_;
  assign new_n_n419_ = ~new_no35_;
  assign new_n_n386_ = ~new_ns1_;
  assign new_n_n375_ = ~new_nf34_;
  assign new_n_n320_ = ~new_nq32_;
  assign new_n_n309_ = ~new_nx31_;
  assign new_n_n287_ = ~new_nb30_;
  assign new_n_n276_ = ~new_nt29_;
  assign new_n_n221_ = ~new_nu24_;
  assign new_n_n210_ = ~new_na24_;
  assign new_n_n199_ = ~new_nq21_;
  assign new_n_n188_ = ~new_nb22_;
  assign new_n_n177_ = ~new_nc21_;
  assign new_n_n123_ = ~new_nc54_;
  assign new_n_n112_ = ~new_nv48_;
  assign new_n_n101_ = ~new_nt46_;
  assign new_n_n90_ = ~new_na45_;
  assign new_nb6_ = ~new_nj54_;
  assign new_ne6_ = new_n_n8_ & new_n_n2_;
  assign new_nv7_ = new_nb_ | new_n_n43_;
  assign new_nb8_ = new_n_n1387_ | new_n_n1386_ | new_n_n1385_;
  assign new_nl8_ = new_n_n57_ | new_n_n61_;
  assign new_nr8_ = new_n_n67_ & new_ne52_;
  assign new_nw8_ = new_n_n72_ | new_n_n73_;
  assign new_nf9_ = new_nz_ | new_n_n82_;
  assign new_ns9_ = new_nz_ | new_n_n94_;
  assign new_nl16_ = new_nu19_ & new_nv0_;
  assign new_nz16_ = new_n_n1373_ | new_n_n1374_;
  assign new_no17_ = new_n_n1369_ | new_n_n1370_;
  assign new_nv17_ = new_n_n434_ | new_nb17_;
  assign new_nk19_ = new_n_n432_ & new_n_n406_;
  assign new_no21_ = new_n_n1333_ | new_n_n1335_ | new_n_n1334_ | new_n_n1336_;
  assign new_n_n1130_ = new_n_n300_ & new_n_n324_;
  assign new_n_n1125_ = new_n_n305_ & new_n_n324_;
  assign new_ny34_ = new_n_n390_ | new_n_n449_;
  assign new_nh35_ = new_n_n409_ | new_n_n437_;
  assign new_np38_ = new_n_n1073_ | new_n_n1072_ | new_n_n1071_;
  assign new_n_n1068_ = new_n_n489_ & new_n_n488_;
  assign new_np40_ = new_n_n1041_ | new_n_n1040_ | new_n_n1039_;
  assign new_nt40_ = new_nc52_ & new_n_n518_;
  assign new_nr41_ = new_n_n1025_ | new_ni0_;
  assign new_n_n1009_ = new_n_n792_ & new_n_n735_ & new_np41_ & new_n_n760_;
  assign new_n_n1003_ = new_n_n735_ & new_nq42_;
  assign new_n_n985_ = new_nl51_ & new_n_n550_;
  assign new_n_n982_ = new_nz50_ & new_n_n552_;
  assign new_n_n973_ = new_n_n563_ & new_n_n558_;
  assign new_nu43_ = new_n_n967_ | new_n_n966_ | new_n_n965_;
  assign new_n_n952_ = new_n_n575_ & new_n_n734_;
  assign new_n_n945_ = new_n_n594_ & new_n_n576_;
  assign new_n_n939_ = new_n_n580_ & new_n_n790_;
  assign new_n_n932_ = new_n_n594_ & new_n_n582_;
  assign new_n_n929_ = new_n_n584_ & new_n_n760_;
  assign new_n_n924_ = new_n_n586_ & new_n_n792_;
  assign new_nk46_ = new_n_n914_ | new_n_n913_ | new_n_n912_;
  assign new_nv46_ = new_n_n676_ & new_nv50_;
  assign new_na48_ = new_n_n604_ & new_n_n605_;
  assign new_nl48_ = new_n_n894_ | new_n_n895_;
  assign new_ny48_ = new_n_n633_ | new_nz_;
  assign new_nj49_ = new_n_n623_ | new_n_n613_;
  assign new_nt50_ = new_nz_ | new_nm5_ | new_n_n682_ | new_n_n685_;
  assign new_nf51_ = new_ns4_ & new_n_n704_;
  assign new_n_n863_ = new_n_n711_ & new_n_n710_ & new_n_n642_;
  assign new_nz51_ = new_n_n856_ | new_n_n857_;
  assign new_nf52_ = new_n_n855_ | new_n_n650_;
  assign new_n_n852_ = new_n_n655_ & new_nr5_ & new_ns48_;
  assign new_n_n844_ = new_n_n657_ & new_n_n685_ & new_n_n672_;
  assign new_nh53_ = new_n_n663_ | new_n_n662_;
  assign new_nq54_ = new_ne52_ | new_n_n791_;
  assign new_nz54_ = new_n_n704_ | new_n_n779_;
  assign new_ne55_ = new_n_n709_ | new_n_n789_;
  assign new_nn55_ = new_n_n728_ & new_n_n727_ & new_n_n726_;
  assign new_na56_ = new_n_n746_ | new_n_n744_ | new_n_n745_ | new_n_n743_;
  assign new_nj56_ = new_n_n760_ | new_n_n791_;
  assign new_n_n780_ = ~new_nu4_;
  assign new_n_n771_ = ~new_ng56_;
  assign new_n_n766_ = ~new_nm56_;
  assign new_n_n757_ = ~new_nk4_;
  assign new_n_n744_ = ~new_np55_;
  assign new_n_n735_ = ~new_nx3_;
  assign new_n_n681_ = ~new_nw54_;
  assign new_n_n672_ = ~new_nt52_;
  assign new_n_n667_ = ~new_nq53_;
  assign new_n_n646_ = ~new_nm53_;
  assign new_n_n637_ = ~new_nh5_;
  assign new_n_n583_ = ~new_nk45_;
  assign new_n_n574_ = ~new_ns44_;
  assign new_n_n547_ = ~new_nh42_;
  assign new_n_n538_ = ~new_nr41_;
  assign new_n_n484_ = ~new_nd38_;
  assign new_n_n475_ = ~new_nr36_;
  assign new_n_n448_ = ~new_nt2_;
  assign new_n_n409_ = ~new_ni2_;
  assign new_n_n385_ = ~new_nl2_;
  assign new_n_n376_ = ~new_ng34_;
  assign new_n_n319_ = ~new_nr32_;
  assign new_n_n310_ = ~new_no31_;
  assign new_n_n286_ = ~new_na30_;
  assign new_n_n277_ = ~new_nr29_;
  assign new_n_n220_ = ~new_nv24_;
  assign new_n_n211_ = ~new_nz23_;
  assign new_n_n189_ = ~new_nc22_;
  assign new_n_n187_ = ~new_na22_;
  assign new_n_n178_ = ~new_nc_;
  assign new_n_n122_ = ~new_nz51_;
  assign new_n_n113_ = ~new_nj49_;
  assign new_n_n100_ = ~new_ns46_;
  assign new_n_n91_ = ~new_ne45_;
  assign new_nw7_ = new_n_n1390_ | new_n_n1389_ | new_n_n1388_;
  assign new_n_n1385_ = new_n_n50_ & new_nt20_;
  assign new_ni8_ = new_n_n57_ | new_n_n58_;
  assign new_n_n1382_ = new_n_n523_ & new_nj50_;
  assign new_nx8_ = new_n_n72_ | new_n_n74_;
  assign new_ni9_ = new_nz_ | new_n_n85_;
  assign new_np9_ = new_nz_ | new_n_n91_;
  assign new_n_n1379_ = new_n_n127_ & new_n_n356_;
  assign new_nb17_ = new_n_n134_ | new_n_n133_;
  assign new_nm17_ = new_n_n1371_ | new_n_n1372_;
  assign new_n_n1365_ = new_n_n140_ & new_n_n407_;
  assign new_n_n1362_ = new_n_n142_ & new_n_n154_;
  assign new_ns18_ = new_n_n149_ & new_n_n150_;
  assign new_nb21_ = new_n_n362_ | new_nh22_ | new_n_n356_;
  assign new_n_n1178_ = new_n_n265_ & new_n_n413_;
  assign new_nv28_ = new_n_n1174_ | new_n_n1173_ | new_n_n1172_;
  assign new_np31_ = new_n_n310_ | new_n_n366_;
  assign new_n_n1126_ = new_n_n306_ & new_ne19_;
  assign new_nv34_ = new_n_n387_ | new_n_n443_;
  assign new_ng35_ = new_n_n408_ | new_n_n435_;
  assign new_nt38_ = new_n_n1068_ | new_n_n1067_ | new_n_n1066_;
  assign new_n_n1041_ = new_n_n515_ & new_n_n514_;
  assign new_nc41_ = new_n_n1030_ | new_n_n1031_;
  assign new_n_n1026_ = new_n_n790_ & new_n_n759_ & new_n_n734_;
  assign new_nt42_ = new_n_n995_ | new_n_n996_;
  assign new_n_n989_ = new_n_n563_ & new_n_n548_;
  assign new_n_n984_ = new_n_n567_ & new_n_n714_;
  assign new_n_n980_ = new_na4_ & new_n_n554_;
  assign new_np43_ = new_n_n975_ | new_n_n974_ | new_n_n973_;
  assign new_ns43_ = new_n_n568_ & new_n_n561_;
  assign new_n_n951_ = new_nv50_ & new_n_n734_;
  assign new_n_n943_ = new_n_n784_ & new_n_n577_;
  assign new_n_n941_ = new_nj4_ & new_n_n579_;
  assign new_n_n933_ = new_nv50_ & new_n_n735_;
  assign new_n_n928_ = new_nv50_ & new_n_n760_;
  assign new_ng46_ = new_n_n920_ | new_n_n921_;
  assign new_nj46_ = new_n_n915_ | new_n_n916_;
  assign new_nu46_ = new_ny45_ & new_no4_;
  assign new_nb48_ = new_ny50_ & new_ny4_;
  assign new_no48_ = new_n_n892_ | new_n_n893_;
  assign new_nv48_ = new_n_n888_ | new_n_n889_;
  assign new_ni49_ = new_n_n615_ | new_n_n614_ | new_nr49_;
  assign new_nt49_ = new_n_n622_ | new_n_n621_;
  assign new_nc50_ = new_n_n878_ | new_n_n877_ | new_n_n876_;
  assign new_n_n866_ = new_n_n686_ & new_n_n711_ & new_n_n644_;
  assign new_nw51_ = new_nm51_ | new_nz_;
  assign new_n_n855_ = new_n_n651_ & new_n_n652_;
  assign new_n_n851_ = new_n_n672_ & new_nm53_;
  assign new_n_n846_ = new_n_n689_ & new_n_n656_ & new_n_n674_;
  assign new_ng53_ = new_n_n689_ | new_nm53_;
  assign new_nn54_ = new_n_n684_ | new_n_n785_;
  assign new_ny54_ = new_n_n703_ & new_n_n702_ & new_n_n701_;
  assign new_nf55_ = new_n_n710_ | new_n_n791_;
  assign new_nq55_ = new_n_n731_ | new_n_n783_;
  assign new_nx55_ = new_n_n738_ | new_n_n797_;
  assign new_ni56_ = new_n_n759_ | new_n_n789_;
  assign new_n_n783_ = ~new_ns0_;
  assign new_n_n772_ = ~new_nh56_;
  assign new_n_n765_ = ~new_nl56_;
  assign new_n_n754_ = ~new_nt4_;
  assign new_n_n747_ = ~new_ns55_;
  assign new_n_n736_ = ~new_na4_;
  assign new_n_n684_ = ~new_ng4_;
  assign new_n_n673_ = ~new_nc0_;
  assign new_n_n666_ = ~new_nn53_;
  assign new_n_n655_ = ~new_na0_;
  assign new_n_n638_ = ~new_np46_;
  assign new_n_n586_ = ~new_nd46_;
  assign new_n_n575_ = ~new_nv44_;
  assign new_n_n568_ = ~new_ng41_;
  assign new_n_n557_ = ~new_ne43_;
  assign new_n_n487_ = ~new_np38_;
  assign new_n_n476_ = ~new_nn37_;
  assign new_n_n458_ = ~new_nv35_;
  assign new_n_n399_ = ~new_nt34_;
  assign new_n_n388_ = ~new_ny1_;
  assign new_n_n377_ = ~new_nh34_;
  assign new_n_n300_ = ~new_nw30_;
  assign new_n_n289_ = ~new_nn29_;
  assign new_n_n278_ = ~new_nf29_;
  assign new_n_n219_ = ~new_nx24_;
  assign new_n_n201_ = ~new_nt22_;
  assign new_n_n190_ = ~new_nk22_;
  assign new_n_n121_ = ~new_nw51_;
  assign new_n_n110_ = ~new_nq48_;
  assign new_n_n103_ = ~new_no47_;
  assign new_n_n92_ = ~new_np45_;
  assign new_nc6_ = new_n_n8_ & new_n_n0_;
  assign new_n_n1390_ = new_np2_ & new_n_n45_;
  assign new_n_n1386_ = new_n_n50_ & new_ne19_;
  assign new_nj8_ = new_nt20_ & new_n_n59_;
  assign new_n_n1383_ = new_ne52_ & new_n_n66_;
  assign new_ny8_ = new_ne52_ & new_n_n75_;
  assign new_nh9_ = new_n_n676_ & new_n_n84_;
  assign new_nq9_ = new_nz_ | new_n_n92_;
  assign new_ns16_ = new_n_n159_ | new_n_n129_ | new_nb_ | new_n_n128_;
  assign new_n_n1373_ = new_n_n132_ & new_n_n432_;
  assign new_n_n1372_ = new_nm16_ & new_nz0_;
  assign new_n_n1366_ = new_nj17_ & new_nc1_;
  assign new_n_n1361_ = new_n_n142_ & new_nr18_;
  assign new_nr18_ = new_nf1_ | new_n_n148_;
  assign new_n_n1345_ = new_n_n169_ & new_n_n167_ & new_n_n363_;
  assign new_n_n1177_ = new_n_n265_ & new_n_n271_;
  assign new_n_n1175_ = new_n_n440_ & new_ns28_;
  assign new_nr31_ = new_n_n1131_ | new_n_n1130_ | new_n_n1129_;
  assign new_nx31_ = new_n_n1126_ | new_n_n1125_ | new_n_n1124_;
  assign new_nw34_ = new_n_n388_ | new_n_n445_;
  assign new_nf35_ = new_n_n407_ | new_n_n433_;
  assign new_n_n1074_ = new_n_n688_ & new_n_n482_;
  assign new_n_n1036_ = new_n_n521_ & new_n_n519_;
  assign new_n_n1031_ = new_nu3_ & new_ng41_;
  assign new_np41_ = new_n_n1026_ | new_ni0_;
  assign new_n_n996_ = new_ny3_ & new_n_n544_;
  assign new_n_n990_ = new_nz50_ & new_n_n547_;
  assign new_na43_ = new_n_n568_ & new_n_n551_;
  assign new_nl43_ = new_n_n979_ | new_n_n980_;
  assign new_n_n975_ = new_n_n558_ & new_n_n557_;
  assign new_n_n968_ = new_n_n567_ & new_n_n764_;
  assign new_n_n950_ = new_n_n594_ & new_n_n575_;
  assign new_n_n944_ = new_ni4_ & new_ni44_;
  assign new_n_n940_ = new_n_n732_ & new_ni45_;
  assign new_n_n934_ = new_n_n582_ & new_n_n735_;
  assign new_n_n927_ = new_n_n594_ & new_n_n584_;
  assign new_n_n922_ = new_n_n594_ & new_n_n586_;
  assign new_n_n916_ = new_no4_ & new_n_n589_;
  assign new_nt46_ = new_n_n788_ | new_n_n758_ | new_n_n733_;
  assign new_nc48_ = new_n_n683_ | new_n_n705_ | new_n_n730_;
  assign new_n_n894_ = new_n_n607_ & new_n_n705_;
  assign new_n_n889_ = new_ny47_ & new_n_n782_;
  assign new_ng49_ = new_nd5_ | new_n_n612_;
  assign new_nu49_ = new_n_n623_ & new_n_n624_;
  assign new_n_n879_ = new_n_n676_ & new_n_n629_ & new_n_n627_;
  assign new_n_n865_ = new_n_n686_ & new_n_n710_ & new_n_n643_;
  assign new_n_n858_ = new_n_n646_ & new_nj5_;
  assign new_ni52_ = new_n_n653_ | new_ng49_ | new_nu53_;
  assign new_nu52_ = new_n_n848_ | new_n_n850_ | new_n_n849_ | new_n_n851_;
  assign new_ny52_ = new_n_n844_ | new_n_n842_ | new_n_n841_ | new_n_n840_ | new_n_n843_ | new_n_n845_;
  assign new_nf53_ = new_nm52_ | new_nu53_;
  assign new_no54_ = new_np46_ | new_n_n787_;
  assign new_nx54_ = new_n_n700_ | new_n_n698_ | new_n_n699_ | new_n_n697_;
  assign new_ng55_ = new_n_n711_ | new_n_n793_;
  assign new_np55_ = new_n_n730_ | new_n_n781_;
  assign new_ny55_ = new_n_n739_ | new_n_n799_;
  assign new_nh56_ = new_n_n758_ | new_n_n787_;
  assign new_n_n782_ = ~new_nz4_;
  assign new_n_n773_ = ~new_ni56_;
  assign new_n_n764_ = ~new_ns3_;
  assign new_n_n755_ = ~new_ny4_;
  assign new_n_n746_ = ~new_nr55_;
  assign new_n_n737_ = ~new_ng3_;
  assign new_n_n683_ = ~new_nv4_;
  assign new_n_n674_ = ~new_nv52_;
  assign new_n_n665_ = ~new_np53_;
  assign new_n_n656_ = ~new_nj51_;
  assign new_n_n648_ = ~new_nk5_;
  assign new_n_n585_ = ~new_nn45_;
  assign new_n_n576_ = ~new_nz44_;
  assign new_n_n567_ = ~new_nl51_;
  assign new_n_n558_ = ~new_ng43_;
  assign new_n_n486_ = ~new_nr38_;
  assign new_n_n477_ = ~new_nc52_;
  assign new_n_n468_ = ~new_nh37_;
  assign new_n_n389_ = ~new_nr2_;
  assign new_n_n387_ = ~new_nv1_;
  assign new_n_n378_ = ~new_na35_;
  assign new_n_n299_ = ~new_nf31_;
  assign new_n_n290_ = ~new_nz30_;
  assign new_n_n288_ = ~new_nq29_;
  assign new_n_n209_ = ~new_nc24_;
  assign new_n_n200_ = ~new_nd_;
  assign new_n_n191_ = ~new_ni22_;
  assign new_n_n120_ = ~new_nv51_;
  assign new_n_n111_ = ~new_np47_;
  assign new_n_n102_ = ~new_nx46_;
  assign new_n_n93_ = ~new_ns45_;
  assign new_np6_ = new_n_n12_ | new_n_n11_;
  assign new_nc7_ = new_nb_ | new_n_n22_;
  assign new_nn7_ = new_nb_ | new_n_n32_;
  assign new_nb10_ = new_n_n111_ & new_n_n106_;
  assign new_no10_ = new_n_n119_ | new_n_n118_;
  assign new_ng16_ = new_n_n1380_ | new_n_n1381_;
  assign new_n_n1353_ = new_n_n181_ & new_np22_;
  assign new_nd29_ = new_n_n274_ & new_n_n272_;
  assign new_n_n1163_ = new_n_n282_ & new_n_n448_;
  assign new_n_n1121_ = new_n_n311_ & new_ne19_;
  assign new_nr32_ = new_n_n316_ & new_nc3_;
  assign new_ny32_ = new_n_n1111_ | new_n_n1110_ | new_n_n1109_;
  assign new_n_n1105_ = new_n_n325_ & new_n_n324_;
  assign new_no33_ = new_n_n336_ | new_n_n437_;
  assign new_np35_ = new_n_n417_ | new_n_n418_ | new_n_n419_;
  assign new_na36_ = new_n_n446_ | new_n_n445_;
  assign new_n_n1099_ = new_n_n712_ & new_n_n737_;
  assign new_nz36_ = new_n_n686_ | new_nm53_;
  assign new_n_n1088_ = new_n_n737_ & new_n_n468_;
  assign new_n_n1082_ = new_nj50_ & new_n_n474_;
  assign new_nf38_ = new_ne37_ & new_nl3_;
  assign new_n_n1075_ = new_nl3_ & new_nn38_;
  assign new_n_n1058_ = new_no3_ & new_n_n494_;
  assign new_no39_ = new_n_n500_ | new_n_n523_;
  assign new_na40_ = new_n_n738_ | new_no3_ | new_np3_;
  assign new_n_n1044_ = new_n_n520_ & new_nd39_;
  assign new_n_n1037_ = new_n_n764_ & new_nt40_;
  assign new_nx40_ = new_n_n524_ | new_n_n523_;
  assign new_no41_ = new_nu3_ & new_nv3_;
  assign new_ny42_ = new_n_n987_ | new_n_n988_;
  assign new_nj43_ = new_nb4_ & new_na4_ & new_nm42_;
  assign new_n_n976_ = new_n_n567_ & new_n_n739_;
  assign new_n_n969_ = new_nl51_ & new_n_n560_;
  assign new_ny43_ = new_n_n568_ & new_n_n569_;
  assign new_nn44_ = new_n_n591_ | new_n_n684_;
  assign new_ns46_ = new_n_n708_ | new_n_n786_ | new_n_n757_;
  assign new_n_n905_ = new_n_n651_ & new_n_n710_;
  assign new_n_n902_ = new_n_n599_ & new_n_n729_;
  assign new_nr53_ = new_n_n676_ & new_n_n685_;
  assign new_n_n836_ = new_np5_ & new_ny53_ & new_n_n676_;
  assign new_ng54_ = new_n_n823_ | new_n_n822_ | new_n_n825_ | new_n_n824_ | new_n_n821_ | new_n_n820_ | new_n_n826_ | new_n_n819_;
  assign new_n_n817_ = new_n_n711_ & new_n_n686_ & new_n_n677_;
  assign new_nr56_ = new_n_n778_ & new_n_n777_ & new_n_n776_;
  assign new_nc57_ = new_n_n800_ | new_n_n799_;
  assign new_n_n804_ = ~new_ns56_;
  assign new_n_n793_ = ~new_nn0_;
  assign new_n_n727_ = ~new_nb56_;
  assign new_n_n716_ = ~new_ni55_;
  assign new_n_n705_ = ~new_nw4_;
  assign new_n_n694_ = ~new_nl54_;
  assign new_n_n678_ = ~new_nx53_;
  assign new_n_n618_ = ~new_nc5_;
  assign new_n_n607_ = ~new_nf48_;
  assign new_n_n596_ = ~new_ny50_;
  assign new_n_n580_ = ~new_no45_;
  assign new_n_n569_ = ~new_nu43_;
  assign new_n_n508_ = ~new_na40_;
  assign new_n_n497_ = ~new_ne38_;
  assign new_n_n481_ = ~new_ne37_;
  assign new_n_n470_ = ~new_nn36_;
  assign new_n_n459_ = ~new_nw35_;
  assign new_n_n398_ = ~new_ns34_;
  assign new_n_n382_ = ~new_nb1_;
  assign new_n_n371_ = ~new_nb34_;
  assign new_n_n360_ = ~new_nk2_;
  assign new_n_n349_ = ~new_np33_;
  assign new_n_n283_ = ~new_ng29_;
  assign new_n_n272_ = ~new_nr22_;
  assign new_n_n261_ = ~new_nc28_;
  assign new_n_n250_ = ~new_nu26_;
  assign new_n_n239_ = ~new_nj25_;
  assign new_n_n184_ = ~new_nt21_;
  assign new_n_n174_ = ~new_ns18_;
  assign new_n_n163_ = ~new_nj1_;
  assign new_n_n152_ = ~new_ny19_;
  assign new_n_n141_ = ~new_nb17_;
  assign new_n_n130_ = ~new_nl16_;
  assign new_nx5_ = ~new_nr56_;
  assign new_no6_ = new_n_n10_ | new_n_n143_;
  assign new_nd7_ = new_nb_ | new_n_n23_;
  assign new_nm7_ = new_nb_ | new_n_n31_;
  assign new_no9_ = new_nz_ | new_n_n90_;
  assign new_na10_ = new_n_n111_ & new_n_n105_;
  assign new_nq10_ = new_n_n121_ & new_n_n120_;
  assign new_nf16_ = new_nn6_ | new_ng1_;
  assign new_n_n1356_ = new_no28_ & new_n_n163_;
  assign new_ne29_ = new_n_n1167_ | new_n_n1168_;
  assign new_nn29_ = new_n_n1163_ | new_nj_;
  assign new_n_n1120_ = new_n_n310_ & new_n_n324_;
  assign new_nq32_ = new_n_n391_ & new_n_n315_;
  assign new_n_n1111_ = new_n_n320_ & new_ne19_;
  assign new_n_n1106_ = new_n_n326_ & new_ne19_;
  assign new_ny33_ = new_n_n352_ | new_n_n350_ | new_n_n351_ | new_n_n349_;
  assign new_nq35_ = new_n_n423_ | new_n_n421_ | new_n_n422_ | new_n_n420_;
  assign new_nz35_ = new_n_n444_ | new_n_n443_;
  assign new_no36_ = new_n_n466_ & new_n_n464_;
  assign new_ns36_ = new_n_n466_ & new_n_n467_;
  assign new_nh37_ = new_nc52_ & new_n_n469_;
  assign new_nn37_ = new_n_n1081_ | new_n_n1082_;
  assign new_ng38_ = new_nk3_ & new_ne37_;
  assign new_nm38_ = new_n_n1074_ | new_n_n1075_;
  assign new_nb39_ = new_nq3_ | new_n_n502_;
  assign new_nq39_ = new_nc52_ & new_n_n501_;
  assign new_nw39_ = new_nc52_ & new_n_n506_;
  assign new_nm40_ = new_n_n1042_ | new_n_n1043_;
  assign new_n_n1038_ = new_ns3_ & new_n_n516_;
  assign new_nz40_ = new_nc52_ & new_n_n525_;
  assign new_nm41_ = new_n_n759_ & new_n_n734_;
  assign new_n_n988_ = new_nz3_ & new_n_n549_;
  assign new_nh43_ = new_nk42_ & new_n_n736_ & new_n_n761_;
  assign new_nn43_ = new_n_n568_ & new_n_n556_;
  assign new_n_n970_ = new_n_n560_ & new_n_n764_;
  assign new_ne44_ = new_nj0_ | new_n_n686_;
  assign new_n_n955_ = new_n_n756_ & new_n_n571_;
  assign new_n_n917_ = new_n_n594_ & new_n_n588_;
  assign new_ng47_ = new_n_n780_ | new_n_n729_ | new_n_n754_ | new_n_n704_;
  assign new_n_n903_ = new_ni47_ & new_ns4_;
  assign new_ns53_ = new_nn5_ | new_n_n671_;
  assign new_nc54_ = new_n_n836_ | new_n_n835_ | new_n_n834_;
  assign new_n_n826_ = new_n_n711_ & new_n_n686_ & new_n_n710_;
  assign new_n_n818_ = new_n_n711_ & new_n_n710_ & new_nw53_;
  assign new_ns56_ = new_n_n780_ | new_n_n779_;
  assign new_nb57_ = new_n_n798_ | new_n_n797_;
  assign new_n_n803_ = ~new_nc57_;
  assign new_n_n794_ = ~new_nc4_;
  assign new_n_n726_ = ~new_nz55_;
  assign new_n_n717_ = ~new_nj55_;
  assign new_n_n704_ = ~new_nr4_;
  assign new_n_n695_ = ~new_nm54_;
  assign new_n_n668_ = ~new_nr53_;
  assign new_n_n628_ = ~new_ng5_;
  assign new_n_n606_ = ~new_nj47_;
  assign new_n_n597_ = ~new_ni52_;
  assign new_n_n579_ = ~new_ni45_;
  assign new_n_n570_ = ~new_ne44_;
  assign new_n_n507_ = ~new_ne40_;
  assign new_n_n498_ = ~new_ng38_;
  assign new_n_n480_ = ~new_nb37_;
  assign new_n_n471_ = ~new_nq36_;
  assign new_n_n449_ = ~new_nn_;
  assign new_n_n408_ = ~new_nd2_;
  assign new_n_n381_ = ~new_nw0_;
  assign new_n_n372_ = ~new_nc34_;
  assign new_n_n359_ = ~new_nf2_;
  assign new_n_n350_ = ~new_nq33_;
  assign new_n_n282_ = ~new_ne29_;
  assign new_n_n273_ = ~new_nd29_;
  assign new_n_n260_ = ~new_nm27_;
  assign new_n_n251_ = ~new_ny26_;
  assign new_n_n229_ = ~new_np25_;
  assign new_n_n183_ = ~new_nd22_;
  assign new_n_n175_ = ~new_nq20_;
  assign new_n_n162_ = ~new_no1_;
  assign new_n_n153_ = ~new_nz19_;
  assign new_n_n140_ = ~new_nj17_;
  assign new_n_n131_ = ~new_no16_;
  assign new_ny5_ = ~new_nc56_;
  assign new_ns6_ = new_n_n268_ & new_nf22_;
  assign new_na7_ = new_n_n268_ & new_n_n20_;
  assign new_nl7_ = new_nb_ | new_n_n30_;
  assign new_ne9_ = new_nz_ | new_n_n81_;
  assign new_nd10_ = new_n_n111_ & new_n_n108_;
  assign new_nm10_ = new_nf50_ & new_n_n116_;
  assign new_nb16_ = new_n_n163_ | new_no28_;
  assign new_nt29_ = new_nr20_ & new_n_n277_;
  assign new_n_n1151_ = new_n_n283_ & new_n_n324_;
  assign new_n_n1119_ = new_n_n310_ & new_n_n311_;
  assign new_nt32_ = new_nd3_ & new_nc3_ & new_n_n316_;
  assign new_n_n1112_ = new_n_n391_ & new_n_n317_;
  assign new_ne33_ = new_n_n1106_ | new_n_n1105_ | new_n_n1104_;
  assign new_ni34_ = new_n_n364_ | new_n_n447_;
  assign new_nr35_ = new_n_n427_ | new_n_n425_ | new_n_n426_ | new_n_n424_;
  assign new_nc36_ = new_n_n450_ | new_n_n449_;
  assign new_n_n1100_ = new_n_n712_ & new_n_n477_;
  assign new_n_n1094_ = new_n_n465_ & new_n_n471_;
  assign new_nj37_ = new_n_n1087_ | new_n_n1086_ | new_n_n1085_;
  assign new_no37_ = new_n_n477_ | new_n_n476_;
  assign new_nd38_ = new_n_n688_ & new_nb37_;
  assign new_n_n1076_ = new_n_n520_ & new_n_n481_;
  assign new_nc39_ = new_n_n1062_ | new_nh0_;
  assign new_ni39_ = new_n_n495_ | new_n_n523_;
  assign new_nu39_ = new_n_n505_ | new_n_n523_;
  assign new_n_n1043_ = new_nr3_ & new_nn40_;
  assign new_ns40_ = new_nj50_ | new_ne52_;
  assign new_n_n1033_ = new_nt3_ & new_n_n522_;
  assign new_ng41_ = new_n_n527_ & new_n_n528_;
  assign new_n_n1020_ = new_n_n530_ & new_n_n713_;
  assign new_nz41_ = new_n_n1012_ | new_n_n1011_ | new_n_n1010_;
  assign new_n_n987_ = new_n_n792_ & new_na43_;
  assign new_n_n983_ = new_n_n553_ & new_n_n552_;
  assign new_n_n978_ = new_n_n555_ & new_n_n739_;
  assign new_nr43_ = new_n_n970_ | new_n_n969_ | new_n_n968_;
  assign new_n_n961_ = new_nl51_ & new_n_n566_;
  assign new_n_n956_ = new_nf4_ & new_ng44_;
  assign new_ne46_ = new_n_n924_ | new_n_n923_ | new_n_n922_;
  assign new_nd47_ = new_n_n905_ | new_n_n906_;
  assign new_nr47_ = new_n_n902_ | new_n_n903_;
  assign new_nu53_ = new_n_n676_ & new_ns53_;
  assign new_n_n834_ = new_nq5_ & new_ny53_ & new_n_n676_;
  assign new_n_n828_ = new_n_n686_ & new_n_n710_ & new_n_n678_;
  assign new_nh54_ = new_n_n816_ | new_n_n815_ | new_n_n818_ | new_n_n817_ | new_n_n814_ | new_n_n813_ | new_n_n826_ | new_n_n812_;
  assign new_nr54_ = new_n_n686_ | new_n_n793_;
  assign new_nt56_ = new_n_n782_ | new_n_n781_;
  assign new_ne57_ = new_n_n807_ | new_n_n805_ | new_n_n806_ | new_n_n804_;
  assign new_n_n806_ = ~new_nu56_;
  assign new_n_n795_ = ~new_nm0_;
  assign new_n_n779_ = ~new_nu0_;
  assign new_n_n768_ = ~new_nd56_;
  assign new_n_n725_ = ~new_ng55_;
  assign new_n_n714_ = ~new_nq3_;
  assign new_n_n707_ = ~new_nh4_;
  assign new_n_n696_ = ~new_nn54_;
  assign new_n_n680_ = ~new_nx54_;
  assign new_n_n669_ = ~new_nl52_;
  assign new_n_n627_ = ~new_nz49_;
  assign new_n_n616_ = ~new_nb49_;
  assign new_n_n598_ = ~new_nj52_;
  assign new_n_n582_ = ~new_nr45_;
  assign new_n_n571_ = ~new_ng44_;
  assign new_n_n528_ = ~new_nk52_;
  assign new_n_n517_ = ~new_nq40_;
  assign new_n_n483_ = ~new_nl38_;
  assign new_n_n472_ = ~new_nl37_;
  assign new_n_n439_ = ~new_ns_;
  assign new_n_n418_ = ~new_nn35_;
  assign new_n_n384_ = ~new_nh2_;
  assign new_n_n373_ = ~new_nd34_;
  assign new_n_n340_ = ~new_nw2_;
  assign new_n_n329_ = ~new_nf33_;
  assign new_n_n285_ = ~new_nr20_;
  assign new_n_n274_ = ~new_nj_;
  assign new_n_n259_ = ~new_nt27_;
  assign new_n_n241_ = ~new_nk20_;
  assign new_n_n230_ = ~new_nn25_;
  assign new_n_n186_ = ~new_no21_;
  assign new_nv6_ = ~new_np22_;
  assign new_n_n161_ = ~new_ni_;
  assign new_n_n150_ = ~new_nn6_;
  assign new_n_n143_ = ~new_nl18_;
  assign new_n_n132_ = ~new_nq16_;
  assign new_nz5_ = ~new_nn55_;
  assign new_nq6_ = new_n_n14_ | new_n_n13_;
  assign new_nb7_ = new_n_n268_ & new_n_n21_;
  assign new_nk7_ = new_nb_ | new_n_n29_;
  assign new_nu8_ = new_ne52_ & new_n_n70_;
  assign new_nc10_ = new_n_n111_ & new_n_n107_;
  assign new_nn10_ = new_n_n676_ & new_n_n117_;
  assign new_ny10_ = new_n_n126_ & new_nc54_;
  assign new_nv29_ = new_n_n1157_ | new_n_n1156_ | new_n_n1155_;
  assign new_n_n1152_ = new_n_n282_ & new_ne19_;
  assign new_ne32_ = new_n_n1117_ | new_n_n1118_;
  assign new_ns32_ = new_n_n315_ & new_n_n391_ & new_n_n416_;
  assign new_nw32_ = new_nr20_ & new_n_n318_;
  assign new_nc33_ = new_nr20_ & new_n_n323_;
  assign new_ns34_ = new_n_n384_ | new_n_n437_;
  assign new_ns35_ = new_n_n430_ & new_n_n429_ & new_n_n428_;
  assign new_nb36_ = new_n_n448_ | new_n_n447_;
  assign new_nn36_ = new_n_n1099_ | new_ns36_;
  assign new_n_n1095_ = new_n_n465_ & new_n_n762_;
  assign new_n_n1087_ = new_n_n471_ & new_n_n470_;
  assign new_n_n1081_ = new_n_n520_ & new_n_n475_;
  assign new_ne38_ = new_nj3_ & new_nb37_;
  assign new_n_n1077_ = new_nj50_ & new_n_n480_;
  assign new_n_n1062_ = new_ng38_ & new_np3_;
  assign new_n_n1057_ = new_n_n763_ & new_nk39_;
  assign new_n_n1052_ = new_n_n798_ & new_nq39_;
  assign new_n_n1042_ = new_n_n739_ & new_n_n512_;
  assign new_nr40_ = new_n_n517_ | new_n_n523_;
  assign new_n_n1032_ = new_n_n800_ & new_nz40_;
  assign new_n_n1027_ = new_n_n567_ & new_n_n688_;
  assign new_n_n1019_ = new_nl51_ & new_n_n530_;
  assign new_n_n1013_ = new_n_n790_ & new_na42_;
  assign new_nz42_ = new_n_n986_ | new_n_n985_ | new_n_n984_;
  assign new_nk43_ = new_n_n983_ | new_n_n982_ | new_n_n981_;
  assign new_n_n977_ = new_nl51_ & new_n_n555_;
  assign new_n_n971_ = new_n_n761_ & new_ns43_;
  assign new_n_n960_ = new_n_n567_ & new_n_n800_;
  assign new_nl44_ = new_n_n955_ | new_n_n956_;
  assign new_n_n930_ = new_n_n786_ & new_nk45_;
  assign new_n_n906_ = new_n_n651_ & new_nm53_;
  assign new_np47_ = new_n_n633_ | new_n_n598_ | new_nz_ | new_n_n597_;
  assign new_nv53_ = new_n_n709_ & new_n_n682_;
  assign new_n_n835_ = new_nr5_ & new_ny53_ & new_n_n676_;
  assign new_n_n827_ = new_n_n686_ & new_nw53_ & new_n_n678_;
  assign new_n_n819_ = new_n_n710_ & new_nw53_ & new_n_n678_;
  assign new_nb55_ = new_n_n706_ | new_n_n783_;
  assign new_nu56_ = new_n_n784_ | new_n_n783_;
  assign new_nd57_ = new_n_n801_ | new_n_n802_ | new_n_n803_;
  assign new_n_n805_ = ~new_nt56_;
  assign new_n_n796_ = ~new_ni3_;
  assign new_n_n778_ = ~new_ne57_;
  assign new_n_n769_ = ~new_ne56_;
  assign new_n_n724_ = ~new_nf55_;
  assign new_n_n715_ = ~new_nh55_;
  assign new_n_n706_ = ~new_nd4_;
  assign new_n_n697_ = ~new_no54_;
  assign new_n_n679_ = ~new_nv54_;
  assign new_n_n670_ = ~new_no53_;
  assign new_n_n626_ = ~new_no10_;
  assign new_n_n617_ = ~new_na5_;
  assign new_n_n608_ = ~new_ni48_;
  assign new_n_n581_ = ~new_ng45_;
  assign new_n_n572_ = ~new_nj0_;
  assign new_n_n527_ = ~new_nf0_;
  assign new_n_n518_ = ~new_np40_;
  assign new_n_n482_ = ~new_nn38_;
  assign new_n_n473_ = ~new_nj37_;
  assign new_n_n429_ = ~new_ng36_;
  assign new_n_n428_ = ~new_ne36_;
  assign new_n_n383_ = ~new_nc2_;
  assign new_n_n374_ = ~new_ne34_;
  assign new_n_n339_ = ~new_nm21_;
  assign new_n_n330_ = ~new_ne33_;
  assign new_n_n284_ = ~new_nz29_;
  assign new_n_n275_ = ~new_ns22_;
  assign new_n_n249_ = ~new_ns26_;
  assign new_n_n240_ = ~new_na26_;
  assign new_n_n231_ = ~new_nm25_;
  assign new_n_n185_ = ~new_nr21_;
  assign new_n_n176_ = ~new_nh_;
  assign new_n_n160_ = ~new_ng16_;
  assign new_n_n151_ = ~new_nw18_;
  assign new_n_n142_ = ~new_nb18_;
  assign new_n_n133_ = ~new_nd17_;
  assign new_na6_ = ~new_ny54_;
  assign new_nj6_ = new_n_n8_ & new_n_n7_;
  assign new_ny6_ = new_n_n18_ & new_nz22_;
  assign new_nj7_ = new_nb_ | new_n_n28_;
  assign new_nn8_ = new_ne52_ & new_n_n63_;
  assign new_nk10_ = new_n_n113_ | new_n_n612_;
  assign new_nx10_ = new_n_n125_ & new_nc54_;
  assign new_np30_ = new_n_n340_ & new_nn29_;
  assign new_n_n1146_ = new_n_n288_ & new_n_n289_;
  assign new_n_n1118_ = new_nb3_ & new_n_n312_;
  assign new_nk33_ = new_n_n333_ & new_n_n332_ & new_n_n331_;
  assign new_nv33_ = new_n_n341_ | new_n_n451_;
  assign new_ng34_ = new_n_n362_ | new_n_n443_;
  assign new_nr34_ = new_n_n383_ | new_n_n435_;
  assign new_nt35_ = new_n_n432_ | new_n_n431_;
  assign new_ne36_ = new_n_n453_ | new_n_n454_ | new_n_n455_;
  assign new_n_n1097_ = new_n_n465_ & new_n_n470_;
  assign new_ne37_ = new_n_n1092_ | new_nh0_;
  assign new_n_n1091_ = new_nj50_ & new_nf3_;
  assign new_n_n1084_ = new_nh3_ & new_nl37_;
  assign new_nt37_ = new_no3_ | new_nm3_ | new_nn3_ | new_nl3_;
  assign new_n_n1078_ = new_n_n481_ & new_n_n480_;
  assign new_nr38_ = new_nc52_ & new_n_n487_;
  assign new_nd39_ = new_n_n503_ | new_n_n714_;
  assign new_nm39_ = new_n_n1056_ | new_n_n1055_ | new_n_n1054_;
  assign new_n_n1050_ = new_nj50_ & new_n_n502_;
  assign new_nh40_ = new_n_n507_ & new_n_n508_;
  assign new_n_n1040_ = new_nj50_ & new_n_n514_;
  assign new_n_n1034_ = new_n_n520_ & new_n_n521_;
  assign new_n_n1028_ = new_nl51_ & new_n_n526_;
  assign new_n_n1021_ = new_n_n759_ & new_nv41_;
  assign new_n_n1014_ = new_nw3_ & new_n_n534_;
  assign new_n_n1012_ = new_n_n535_ & new_n_n738_;
  assign new_n_n1008_ = new_nz3_ & new_nx3_ & new_nr41_ & new_ny3_;
  assign new_n_n1000_ = new_n_n567_ & new_n_n763_;
  assign new_n_n993_ = new_nl51_ & new_n_n545_;
  assign new_nw43_ = new_n_n962_ | new_n_n961_ | new_n_n960_;
  assign new_n_n957_ = new_n_n731_ & new_n_n706_;
  assign new_n_n937_ = new_n_n594_ & new_n_n580_;
  assign new_n_n907_ = new_n_n594_ & new_n_n595_;
  assign new_n_n904_ = new_n_n596_ & new_n_n704_;
  assign new_nw53_ = new_n_n672_ & new_n_n673_;
  assign new_n_n833_ = new_n_n711_ & new_n_n686_ & new_nw53_;
  assign new_n_n823_ = new_n_n711_ & new_n_n686_ & new_nx53_;
  assign new_n_n813_ = new_n_n711_ & new_n_n686_ & new_n_n678_;
  assign new_nl55_ = new_n_n721_ | new_n_n719_ | new_n_n720_ | new_n_n718_;
  assign new_nv56_ = new_n_n786_ | new_n_n785_;
  assign new_n_n811_ = ~new_nz56_;
  assign new_n_n800_ = ~new_nt3_;
  assign new_n_n789_ = ~new_np0_;
  assign new_n_n759_ = ~new_nv3_;
  assign new_n_n748_ = ~new_nt55_;
  assign new_n_n723_ = ~new_ne55_;
  assign new_n_n712_ = ~new_nf3_;
  assign new_n_n701_ = ~new_nk55_;
  assign new_n_n690_ = ~new_ns54_;
  assign new_n_n660_ = ~new_nw52_;
  assign new_n_n650_ = ~new_nk51_;
  assign new_n_n639_ = ~new_ng51_;
  assign new_n_n625_ = ~new_nr49_;
  assign new_n_n614_ = ~new_nv49_;
  assign new_n_n603_ = ~new_nb48_;
  assign new_n_n592_ = ~new_np4_;
  assign new_n_n562_ = ~new_nh43_;
  assign new_n_n551_ = ~new_nx42_;
  assign new_n_n540_ = ~new_no42_;
  assign new_n_n529_ = ~new_nv41_;
  assign new_n_n526_ = ~new_nc41_;
  assign new_n_n515_ = ~new_ng40_;
  assign new_n_n504_ = ~new_nw39_;
  assign new_n_n493_ = ~new_nk38_;
  assign new_n_n463_ = ~new_na36_;
  assign new_n_n452_ = ~new_ne3_;
  assign new_n_n441_ = ~new_nr_;
  assign new_n_n430_ = ~new_nf36_;
  assign new_n_n427_ = ~new_nl35_;
  assign new_n_n416_ = ~new_nd3_;
  assign new_n_n405_ = ~new_nq35_;
  assign new_n_n394_ = ~new_nz34_;
  assign new_n_n364_ = ~new_nq2_;
  assign new_n_n353_ = ~new_nl34_;
  assign new_n_n342_ = ~new_nt33_;
  assign new_n_n331_ = ~new_nw33_;
  assign new_n_n328_ = ~new_nt20_;
  assign new_n_n317_ = ~new_nw32_;
  assign new_n_n306_ = ~new_nq30_;
  assign new_n_n295_ = ~new_nb31_;
  assign new_n_n279_ = ~new_nc29_;
  assign new_n_n265_ = ~new_ni28_;
  assign new_n_n254_ = ~new_nh27_;
  assign new_n_n243_ = ~new_nd21_;
  assign new_n_n232_ = ~new_ni25_;
  assign new_n_n218_ = ~new_ng24_;
  assign new_n_n207_ = ~new_nq23_;
  assign new_n_n196_ = ~new_nq22_;
  assign new_n_n180_ = ~new_nl32_;
  assign new_n_n170_ = ~new_nn20_;
  assign new_n_n167_ = ~new_nm19_;
  assign new_n_n156_ = ~new_nu18_;
  assign new_n_n145_ = ~new_ny18_;
  assign new_n_n134_ = ~new_ne17_;
  assign new_n_n109_ = ~new_no48_;
  assign new_n_n98_ = ~new_nv46_;
  assign new_nt5_ = ~new_nd35_;
  assign new_ni6_ = new_n_n8_ & new_n_n6_;
  assign new_nz6_ = new_n_n268_ & new_n_n19_;
  assign new_ni7_ = new_nb_ | new_n_n358_;
  assign new_nd8_ = new_nt20_ & new_n_n52_;
  assign new_nl10_ = new_n_n115_ | new_n_n114_;
  assign new_nw10_ = new_n_n124_ | new_n_n123_;
  assign new_nq30_ = new_nu2_ & new_nn29_;
  assign new_n_n1147_ = new_n_n288_ & new_n_n324_;
  assign new_nu32_ = new_n_n1116_ | new_n_n1115_ | new_n_n1114_;
  assign new_nl33_ = new_n_n334_ | new_n_n431_;
  assign new_nu33_ = new_n_n340_ | new_n_n449_;
  assign new_nh34_ = new_n_n363_ | new_n_n445_;
  assign new_nq34_ = new_n_n382_ | new_n_n433_;
  assign new_nu35_ = new_n_n434_ | new_n_n433_;
  assign new_nd36_ = new_n_n452_ | new_n_n451_;
  assign new_nq36_ = new_n_n1096_ | new_ns36_;
  assign new_n_n1093_ = new_n_n474_ & new_n_n796_;
  assign new_n_n1090_ = new_n_n520_ & new_n_n712_;
  assign new_nk37_ = new_n_n1083_ | new_n_n1084_;
  assign new_ny37_ = new_n_n763_ | new_n_n713_ | new_n_n738_ | new_n_n688_;
  assign new_nl38_ = new_n_n1078_ | new_n_n1077_ | new_n_n1076_;
  assign new_n_n1063_ = new_ne38_ & new_n_n798_;
  assign new_ne39_ = new_n_n798_ | new_n_n714_;
  assign new_nk39_ = new_nc52_ & new_n_n496_;
  assign new_n_n1049_ = new_n_n520_ & new_n_n503_;
  assign new_ng40_ = new_n_n510_ & new_nr3_;
  assign new_nl40_ = new_n_n1046_ | new_n_n1045_ | new_n_n1044_;
  assign new_nw40_ = new_n_n1032_ | new_n_n1033_;
  assign new_n_n1029_ = new_n_n526_ & new_n_n688_;
  assign new_nu41_ = new_n_n1020_ | new_n_n1019_ | new_n_n1018_;
  assign new_ny41_ = new_n_n1013_ | new_n_n1014_;
  assign new_n_n1011_ = new_nl51_ & new_n_n535_;
  assign new_nm42_ = new_n_n1008_ | new_ni0_;
  assign new_nq42_ = new_n_n568_ & new_n_n541_;
  assign new_n_n994_ = new_n_n545_ & new_n_n798_;
  assign new_n_n962_ = new_n_n566_ & new_n_n800_;
  assign new_n_n958_ = new_ne4_ & new_nd4_;
  assign new_ni45_ = new_n_n578_ & new_nh4_;
  assign new_nc47_ = new_nj10_ | new_nc5_;
  assign new_ni47_ = new_ny50_ & new_nr4_;
  assign new_nx53_ = new_n_n674_ & new_n_n675_;
  assign new_nf54_ = new_n_n831_ | new_n_n830_ | new_n_n833_ | new_n_n832_ | new_n_n829_ | new_n_n828_ | new_n_n826_ | new_n_n827_;
  assign new_n_n822_ = new_n_n686_ & new_nw53_ & new_nx53_;
  assign new_n_n814_ = new_n_n686_ & new_n_n677_ & new_nx53_;
  assign new_nv55_ = new_n_n736_ | new_n_n793_;
  assign new_nw56_ = new_n_n788_ | new_n_n787_;
  assign new_nf57_ = new_n_n811_ | new_n_n809_ | new_n_n810_ | new_n_n808_;
  assign new_n_n799_ = ~new_nk0_;
  assign new_n_n790_ = ~new_nw3_;
  assign new_n_n758_ = ~new_no4_;
  assign new_n_n749_ = ~new_nu55_;
  assign new_n_n722_ = ~new_nd55_;
  assign new_n_n713_ = ~new_nm3_;
  assign new_n_n700_ = ~new_nr54_;
  assign new_n_n691_ = ~new_nt54_;
  assign new_n_n659_ = ~new_ny52_;
  assign new_n_n651_ = ~new_nc47_;
  assign new_n_n629_ = ~new_nx49_;
  assign new_n_n624_ = ~new_ne5_;
  assign new_n_n615_ = ~new_nu49_;
  assign new_n_n602_ = ~new_na48_;
  assign new_n_n593_ = ~new_nu46_;
  assign new_n_n561_ = ~new_np43_;
  assign new_n_n552_ = ~new_nk42_;
  assign new_n_n539_ = ~new_nq42_;
  assign new_n_n530_ = ~new_nt41_;
  assign new_n_n525_ = ~new_nv40_;
  assign new_n_n516_ = ~new_nt40_;
  assign new_n_n503_ = ~new_nc39_;
  assign new_n_n494_ = ~new_nk39_;
  assign new_n_n462_ = ~new_nz35_;
  assign new_n_n453_ = ~new_nb36_;
  assign new_n_n440_ = ~new_no2_;
  assign new_n_n431_ = ~new_nw_;
  assign new_n_n426_ = ~new_nk35_;
  assign new_n_n417_ = ~new_nm35_;
  assign new_n_n404_ = ~new_nr35_;
  assign new_n_n395_ = ~new_np34_;
  assign new_n_n363_ = ~new_np1_;
  assign new_n_n354_ = ~new_nn34_;
  assign new_n_n341_ = ~new_np21_;
  assign new_n_n332_ = ~new_ny33_;
  assign new_n_n327_ = ~new_ni33_;
  assign new_n_n318_ = ~new_nu32_;
  assign new_n_n305_ = ~new_ns30_;
  assign new_n_n296_ = ~new_nu30_;
  assign new_n_n269_ = ~new_ns28_;
  assign new_n_n264_ = ~new_nx27_;
  assign new_n_n255_ = ~new_nn27_;
  assign new_n_n242_ = ~new_nx25_;
  assign new_n_n233_ = ~new_ng25_;
  assign new_n_n228_ = ~new_nm24_;
  assign new_n_n206_ = ~new_nu23_;
  assign new_n_n197_ = ~new_nn21_;
  assign new_n_n179_ = ~new_np32_;
  assign new_n_n171_ = ~new_ni20_;
  assign new_n_n166_ = ~new_ne20_;
  assign new_n_n157_ = ~new_ng20_;
  assign new_n_n144_ = ~new_nc18_;
  assign new_n_n135_ = ~new_nf17_;
  assign new_n_n108_ = ~new_nl48_;
  assign new_n_n99_ = ~new_nr46_;
  assign new_nu5_ = ~new_no34_;
  assign new_nn6_ = new_ni1_ | new_n_n11_;
  assign new_nw6_ = new_n_n16_ | new_n_n15_;
  assign new_nh7_ = new_nb_ | new_n_n27_;
  assign new_n_n1388_ = new_n_n44_ & new_n_n45_;
  assign new_nz9_ = new_n_n111_ & new_n_n104_;
  assign new_nc31_ = new_n_n1139_ | new_n_n1140_;
  assign new_nh31_ = new_nr20_ & new_n_n299_;
  assign new_n_n1110_ = new_n_n319_ & new_n_n324_;
  assign new_nm33_ = new_n_n335_ | new_n_n433_;
  assign new_nx33_ = new_n_n348_ | new_n_n346_ | new_n_n347_ | new_n_n345_;
  assign new_ne34_ = new_n_n360_ | new_n_n439_;
  assign new_np34_ = new_n_n381_ | new_n_n431_;
  assign new_nv35_ = new_n_n436_ | new_n_n435_;
  assign new_ng36_ = new_n_n463_ | new_n_n461_ | new_n_n462_ | new_n_n460_;
  assign new_np36_ = new_n_n1097_ | new_n_n1098_;
  assign new_nb37_ = new_n_n1093_ | new_nh0_;
  assign new_ng37_ = new_n_n1088_ | new_n_n1089_;
  assign new_nl37_ = new_nc52_ & new_n_n473_;
  assign new_n_n1079_ = new_n_n796_ & new_n_n478_;
  assign new_nk38_ = new_nn3_ & new_nl3_ & new_ne37_ & new_nm3_;
  assign new_n_n1070_ = new_nm3_ & new_nr38_;
  assign new_nz38_ = new_n_n1063_ | new_nh0_;
  assign new_ng39_ = new_n_n1061_ | new_n_n1060_ | new_n_n1059_;
  assign new_n_n1055_ = new_nj50_ & new_n_n497_;
  assign new_ns39_ = new_n_n1051_ | new_n_n1050_ | new_n_n1049_;
  assign new_nf40_ = new_n_n739_ & new_n_n509_;
  assign new_n_n1046_ = new_nd39_ & new_nb39_;
  assign new_nq40_ = new_n_n1037_ | new_n_n1038_;
  assign new_ne41_ = new_n_n1029_ | new_n_n1028_ | new_n_n1027_;
  assign new_nt41_ = new_n_n1021_ | new_n_n1022_;
  assign new_n_n1015_ = new_n_n563_ & new_n_n533_;
  assign new_n_n1010_ = new_n_n567_ & new_n_n738_;
  assign new_n_n1007_ = new_n_n538_ & new_n_n537_;
  assign new_n_n1002_ = new_n_n540_ & new_n_n763_;
  assign new_nu42_ = new_n_n994_ | new_n_n993_ | new_n_n992_;
  assign new_n_n964_ = new_nc4_ & new_n_n565_;
  assign new_nj44_ = new_n_n957_ | new_n_n958_;
  assign new_n_n949_ = new_nh4_ & new_nn44_;
  assign new_ny53_ = new_n_n839_ | new_n_n838_ | new_n_n837_;
  assign new_n_n831_ = new_n_n711_ & new_n_n710_ & new_nx53_;
  assign new_n_n825_ = new_n_n686_ & new_n_n710_ & new_nw53_;
  assign new_n_n815_ = new_n_n710_ & new_nw53_ & new_nx53_;
  assign new_nf56_ = new_n_n756_ | new_n_n783_;
  assign new_nx56_ = new_n_n790_ | new_n_n789_;
  assign new_n_n809_ = ~new_nx56_;
  assign new_n_n802_ = ~new_nb57_;
  assign new_n_n791_ = ~new_no0_;
  assign new_n_n739_ = ~new_nr3_;
  assign new_n_n728_ = ~new_na56_;
  assign new_n_n721_ = ~new_nc55_;
  assign new_n_n710_ = ~new_nr5_;
  assign new_n_n703_ = ~new_nl55_;
  assign new_n_n692_ = ~new_nu54_;
  assign new_n_n658_ = ~new_ni53_;
  assign new_n_n641_ = ~new_nf51_;
  assign new_n_n630_ = ~new_nf5_;
  assign new_n_n623_ = ~new_nd5_;
  assign new_n_n612_ = ~new_ni49_;
  assign new_n_n605_ = ~new_ng47_;
  assign new_n_n594_ = ~new_nv50_;
  assign new_n_n560_ = ~new_nq43_;
  assign new_n_n549_ = ~new_na43_;
  assign new_n_n542_ = ~new_ne42_;
  assign new_n_n531_ = ~new_ns41_;
  assign new_n_n524_ = ~new_nw40_;
  assign new_n_n513_ = ~new_nl40_;
  assign new_n_n506_ = ~new_ns39_;
  assign new_n_n495_ = ~new_nh39_;
  assign new_n_n479_ = ~new_np37_;
  assign new_n_n461_ = ~new_ny35_;
  assign new_n_n450_ = ~new_na3_;
  assign new_n_n443_ = ~new_nq_;
  assign new_n_n432_ = ~new_ny0_;
  assign new_n_n425_ = ~new_nj35_;
  assign new_n_n414_ = ~new_ns2_;
  assign new_n_n407_ = ~new_nc1_;
  assign new_n_n396_ = ~new_nq34_;
  assign new_n_n380_ = ~new_nb35_;
  assign new_n_n369_ = ~new_nk34_;
  assign new_n_n362_ = ~new_nr1_;
  assign new_n_n351_ = ~new_nr33_;
  assign new_n_n344_ = ~new_nv33_;
  assign new_n_n333_ = ~new_nx33_;
  assign new_n_n326_ = ~new_ns32_;
  assign new_n_n315_ = ~new_nn31_;
  assign new_n_n308_ = ~new_ny31_;
  assign new_n_n297_ = ~new_nt30_;
  assign new_n_n281_ = ~new_nv29_;
  assign new_n_n270_ = ~new_nu28_;
  assign new_n_n263_ = ~new_nf28_;
  assign new_n_n252_ = ~new_nj26_;
  assign new_n_n245_ = ~new_nf26_;
  assign new_n_n234_ = ~new_nu25_;
  assign new_n_n227_ = ~new_no24_;
  assign new_n_n216_ = ~new_np24_;
  assign new_n_n198_ = ~new_ne_;
  assign new_n_n182_ = ~new_nr18_;
  assign new_n_n172_ = ~new_nf16_;
  assign new_n_n165_ = ~new_nf20_;
  assign new_n_n154_ = ~new_nh1_;
  assign new_n_n147_ = ~new_ne18_;
  assign new_n_n136_ = ~new_nj16_;
  assign new_n_n129_ = ~new_nb21_;
  assign new_n_n118_ = ~new_nd51_;
  assign new_nv5_ = ~new_nz33_;
  assign new_nk6_ = new_n_n8_ & new_n_n9_;
  assign new_nx6_ = new_n_n17_ & new_nz22_;
  assign new_ng7_ = new_nb_ | new_n_n26_;
  assign new_np7_ = new_nb_ | new_n_n34_;
  assign new_ny9_ = new_n_n111_ & new_n_n103_;
  assign new_n_n1140_ = new_nx2_ & new_nd31_;
  assign new_n_n1134_ = new_n_n390_ & new_n_n298_;
  assign new_n_n1104_ = new_n_n325_ & new_n_n326_;
  assign new_nn33_ = new_nr20_ | new_n_n435_;
  assign new_nw33_ = new_n_n342_ | new_n_n343_ | new_n_n344_;
  assign new_nf34_ = new_n_n361_ | new_n_n441_;
  assign new_no34_ = new_n_n380_ & new_n_n379_ & new_n_n378_;
  assign new_nw35_ = new_n_n438_ | new_n_n437_;
  assign new_nf36_ = new_n_n459_ | new_n_n457_ | new_n_n458_ | new_n_n456_;
  assign new_n_n1098_ = new_n_n465_ & new_nh3_;
  assign new_na37_ = new_n_n711_ | new_nm53_;
  assign new_n_n1089_ = new_ng3_ & new_nh37_;
  assign new_n_n1083_ = new_n_n762_ & new_n_n472_;
  assign new_nq37_ = new_n_n479_ | new_n_n523_;
  assign new_nj38_ = new_nb37_ & new_n_n713_ & new_n_n738_ & new_n_n688_;
  assign new_n_n1069_ = new_n_n713_ & new_n_n486_;
  assign new_nv38_ = new_nc52_ & new_n_n491_;
  assign new_n_n1061_ = new_n_n493_ & new_n_n492_;
  assign new_n_n1056_ = new_n_n498_ & new_n_n497_;
  assign new_n_n1051_ = new_n_n503_ & new_n_n502_;
  assign new_ne40_ = new_nt3_ | new_nr3_ | new_ns3_ | new_nq3_;
  assign new_n_n1045_ = new_nj50_ & new_nb39_;
  assign new_n_n1039_ = new_n_n520_ & new_n_n515_;
  assign new_n_n1035_ = new_nj50_ & new_n_n519_;
  assign new_n_n1022_ = new_nv3_ & new_n_n529_;
  assign new_n_n1016_ = new_nz50_ & new_n_n532_;
  assign new_na42_ = new_n_n568_ & new_n_n536_;
  assign new_nn42_ = new_n_n1007_ | new_n_n1006_ | new_n_n1005_;
  assign new_n_n1001_ = new_nl51_ & new_n_n540_;
  assign new_n_n995_ = new_n_n760_ & new_nv42_;
  assign new_n_n963_ = new_n_n794_ & new_ny43_;
  assign new_n_n959_ = new_nf4_ & new_ne4_ & new_nd4_;
  assign new_ns44_ = new_n_n711_ & new_n_n572_;
  assign new_n_n839_ = new_n_n686_ & new_n_n711_;
  assign new_n_n832_ = new_n_n686_ & new_n_n710_ & new_n_n677_;
  assign new_n_n824_ = new_n_n711_ & new_n_n710_ & new_n_n677_;
  assign new_n_n816_ = new_n_n686_ & new_n_n710_ & new_nx53_;
  assign new_np56_ = new_n_n771_ | new_n_n769_ | new_n_n770_ | new_n_n768_;
  assign new_ny56_ = new_n_n792_ | new_n_n791_;
  assign new_n_n810_ = ~new_ny56_;
  assign new_n_n801_ = ~new_na57_;
  assign new_n_n792_ = ~new_nz3_;
  assign new_n_n738_ = ~new_nn3_;
  assign new_n_n729_ = ~new_ns4_;
  assign new_n_n720_ = ~new_nb55_;
  assign new_n_n711_ = ~new_np5_;
  assign new_n_n702_ = ~new_nm55_;
  assign new_n_n693_ = ~new_nk54_;
  assign new_n_n649_ = ~new_np51_;
  assign new_n_n640_ = ~new_nm51_;
  assign new_n_n631_ = ~new_ni51_;
  assign new_n_n622_ = ~new_nb51_;
  assign new_n_n613_ = ~new_nz48_;
  assign new_n_n604_ = ~new_nc48_;
  assign new_n_n595_ = ~new_nw46_;
  assign new_n_n559_ = ~new_ns43_;
  assign new_n_n550_ = ~new_ny42_;
  assign new_n_n541_ = ~new_nn42_;
  assign new_n_n532_ = ~new_nm41_;
  assign new_n_n523_ = ~new_ne52_;
  assign new_n_n514_ = ~new_nf40_;
  assign new_n_n505_ = ~new_nt39_;
  assign new_n_n496_ = ~new_ng39_;
  assign new_n_n469_ = ~new_nf37_;
  assign new_n_n460_ = ~new_nx35_;
  assign new_n_n451_ = ~new_nm_;
  assign new_n_n442_ = ~new_nu1_;
  assign new_n_n433_ = ~new_nv_;
  assign new_n_n424_ = ~new_ni35_;
  assign new_n_n415_ = ~new_nz2_;
  assign new_n_n406_ = ~new_nx0_;
  assign new_n_n397_ = ~new_nr34_;
  assign new_n_n379_ = ~new_nc35_;
  assign new_n_n370_ = ~new_na34_;
  assign new_n_n361_ = ~new_nm1_;
  assign new_n_n352_ = ~new_ns33_;
  assign new_n_n343_ = ~new_nu33_;
  assign new_n_n334_ = ~new_nl1_;
  assign new_n_n325_ = ~new_nt32_;
  assign new_n_n316_ = ~new_np31_;
  assign new_n_n307_ = ~new_nb32_;
  assign new_n_n298_ = ~new_nh31_;
  assign new_n_n280_ = ~new_nx29_;
  assign new_n_n271_ = ~new_nq19_;
  assign new_n_n262_ = ~new_na28_;
  assign new_n_n253_ = ~new_no26_;
  assign new_n_n244_ = ~new_nw25_;
  assign new_n_n235_ = ~new_ns25_;
  assign new_n_n226_ = ~new_nz24_;
  assign new_n_n217_ = ~new_ni24_;
  assign new_n_n208_ = ~new_no23_;
  assign new_n_n181_ = ~new_nh20_;
  assign new_n_n173_ = ~new_nj18_;
  assign new_n_n164_ = ~new_no28_;
  assign new_n_n155_ = ~new_ni1_;
  assign new_n_n146_ = ~new_nx18_;
  assign new_n_n137_ = ~new_nm16_;
  assign new_n_n128_ = ~new_na21_;
  assign new_n_n119_ = ~new_nf50_;
  assign new_nw5_ = ~new_nk33_;
  assign new_ni20_ = new_n_n356_ & new_ng19_;
  assign new_n_n1347_ = new_n_n169_ & new_n_n168_ & new_n_n167_;
  assign new_na21_ = new_n_n174_ | new_nj18_ | new_np22_;
  assign new_n_n1302_ = new_n_n363_ & new_n_n338_ & new_n_n201_;
  assign new_n_n1293_ = new_n_n203_ & new_n_n340_;
  assign new_nv23_ = new_n_n1286_ | new_n_n1287_;
  assign new_n_n1280_ = new_n_n207_ & new_n_n208_;
  assign new_nj24_ = new_nr23_ & new_n_n387_ & new_n_n412_;
  assign new_n_n1269_ = new_nv1_ & new_n_n214_;
  assign new_no25_ = new_n_n1243_ | new_n_n1242_ | new_n_n1241_;
  assign new_n_n1236_ = new_n_n413_ & new_nu25_;
  assign new_n_n1229_ = new_na2_ & new_n_n240_;
  assign new_nk26_ = new_n_n1222_ | new_n_n1223_;
  assign new_n_n1219_ = new_ne2_ & new_n_n266_;
  assign new_n_n1211_ = new_n_n251_ & new_n_n411_;
  assign new_n_n1206_ = new_nh2_ & new_n_n254_;
  assign new_n_n1198_ = new_n_n257_ & new_n_n387_;
  assign new_nc28_ = new_n_n1190_ | new_n_n1191_;
  assign new_n_n1174_ = new_nq19_ & new_n_n446_;
  assign new_n_n1167_ = new_n_n273_ & new_n_n279_;
  assign new_nr29_ = new_n_n1160_ | new_n_n1161_;
  assign new_nw29_ = new_n_n1153_ | new_n_n1154_;
  assign new_nc30_ = new_n_n287_ | new_n_n328_;
  assign new_nw30_ = new_ny2_ & new_nw2_ & new_nq29_ & new_nx2_;
  assign new_n_n1142_ = new_n_n292_ & new_n_n324_;
  assign new_n_n1135_ = new_ny2_ & new_nh31_;
  assign new_n_n1109_ = new_n_n319_ & new_n_n320_;
  assign new_n_n1103_ = new_ne3_ & new_n_n327_;
  assign new_nr33_ = new_nt20_ | new_n_n443_;
  assign new_nc34_ = new_n_n358_ | new_n_n435_;
  assign new_nn34_ = new_n_n377_ | new_n_n375_ | new_n_n376_ | new_n_n374_;
  assign new_np37_ = new_n_n1079_ | new_n_n1080_;
  assign new_ni38_ = new_nm3_ & new_nl3_ & new_ne37_;
  assign new_n_n84_ = ~new_nm43_;
  assign new_n_n73_ = ~new_no39_;
  assign new_n_n62_ = ~new_ni36_;
  assign new_n_n51_ = ~new_nk30_;
  assign new_n_n40_ = ~new_np28_;
  assign new_nk20_ = new_n_n1353_ | new_n_n1354_;
  assign new_n_n1348_ = new_n_n362_ & new_n_n168_ & new_n_n167_;
  assign new_nn21_ = new_nl1_ & new_nn1_ & new_n_n268_ & new_nm1_;
  assign new_n_n1301_ = new_n_n338_ & new_n_n362_ & new_nu22_;
  assign new_n_n1294_ = new_n_n241_ & new_n_n340_;
  assign new_n_n1287_ = new_nt1_ & new_n_n204_;
  assign new_n_n1281_ = new_n_n207_ & new_n_n237_;
  assign new_nl24_ = new_nw1_ & new_nv1_ & new_nt23_;
  assign new_nq24_ = new_n_n1268_ | new_n_n1269_;
  assign new_n_n1243_ = new_n_n241_ & new_n_n391_;
  assign new_n_n1237_ = new_nz1_ & new_n_n234_;
  assign new_n_n1228_ = new_n_n446_ & new_na26_;
  assign new_n_n1224_ = new_nd2_ & new_nc2_ & new_nb2_;
  assign new_n_n1218_ = new_n_n336_ & new_nt26_;
  assign new_n_n1212_ = new_nq19_ & new_n_n411_;
  assign new_n_n1205_ = new_n_n384_ & new_nh27_;
  assign new_n_n1199_ = new_nq19_ & new_n_n387_;
  assign new_ng28_ = new_n_n1184_ | new_n_n1183_ | new_n_n1182_;
  assign new_n_n1173_ = new_n_n270_ & new_n_n446_;
  assign new_n_n1168_ = new_n_n273_ & new_ns2_;
  assign new_n_n1161_ = new_ne19_ & new_nq2_;
  assign new_n_n1155_ = new_n_n278_ & new_n_n279_;
  assign new_nd30_ = new_ne19_ | new_nt20_;
  assign new_nv30_ = new_nn29_ & new_n_n365_ & new_n_n390_ & new_n_n340_;
  assign new_n_n1141_ = new_n_n292_ & new_n_n293_;
  assign new_ng31_ = new_n_n1134_ | new_n_n1135_;
  assign new_n_n1116_ = new_nn31_ & new_ne19_;
  assign new_n_n1102_ = new_n_n452_ & new_ni33_;
  assign new_nq33_ = new_n_n337_ | new_n_n441_;
  assign new_nd34_ = new_n_n359_ | new_n_n437_;
  assign new_nm34_ = new_n_n373_ | new_n_n371_ | new_n_n372_ | new_n_n370_;
  assign new_n_n1080_ = new_ni3_ & new_no37_;
  assign new_nh38_ = new_nb37_ & new_n_n688_ & new_n_n713_;
  assign new_n_n85_ = ~new_nr43_;
  assign new_n_n72_ = ~new_ns40_;
  assign new_n_n63_ = ~new_ng37_;
  assign new_n_n50_ = ~new_nf30_;
  assign new_n_n41_ = ~new_nq28_;
  assign new_ng20_ = new_n_n174_ & new_nv6_;
  assign new_nq20_ = new_n_n1344_ | new_n_n1343_ | new_n_n1342_ | new_n_n1341_ | new_n_n1348_ | new_n_n1346_ | new_n_n1345_ | new_n_n1347_ | new_n_n166_;
  assign new_n_n1331_ = new_n_n341_ & new_n_n181_ & new_n_n199_;
  assign new_ne23_ = new_n_n1301_ | new_n_n1300_ | new_n_n1303_ | new_n_n1302_ | new_n_n1299_ | new_n_n1298_ | new_n_n1311_ | new_n_n1297_;
  assign new_ni23_ = new_n_n1294_ | new_n_n1293_ | new_n_n1292_;
  assign new_n_n1286_ = new_n_n411_ & new_nx23_;
  assign new_n_n1279_ = new_nu1_ & new_n_n209_;
  assign new_ng24_ = new_n_n387_ & new_nr23_;
  assign new_n_n1270_ = new_n_n212_ & new_n_n213_;
  assign new_ns25_ = new_n_n1236_ | new_n_n1237_;
  assign new_ny25_ = new_n_n1227_ | new_n_n1226_ | new_n_n1225_;
  assign new_n_n1222_ = new_n_n383_ & new_n_n358_;
  assign new_nt26_ = new_n_n249_ | new_n_n248_;
  assign new_nz26_ = new_n_n1212_ | new_n_n1211_ | new_n_n1210_;
  assign new_no27_ = new_n_n1204_ | new_n_n1203_ | new_n_n1202_;
  assign new_nx27_ = new_nl2_ & new_nk2_ & new_nm27_;
  assign new_n_n1185_ = new_n_n385_ & new_na28_;
  assign new_n_n1172_ = new_n_n270_ & new_n_n271_;
  assign new_n_n1166_ = new_nq2_ & new_nr2_;
  assign new_nq29_ = new_n_n1162_ | new_nj_;
  assign new_n_n1156_ = new_n_n278_ & new_n_n324_;
  assign new_nf30_ = new_nz2_ | new_nx2_ | new_ny2_ | new_nw2_;
  assign new_n_n1148_ = new_n_n289_ & new_ne19_;
  assign new_nb31_ = new_n_n1143_ | new_n_n1142_ | new_n_n1141_;
  assign new_n_n1136_ = new_n_n296_ & new_n_n297_;
  assign new_n_n1117_ = new_n_n366_ & new_nh32_;
  assign new_ng33_ = new_n_n329_ | new_n_n328_;
  assign new_nt33_ = new_n_n339_ | new_n_n447_;
  assign new_na34_ = new_n_n356_ | new_n_n431_;
  assign new_nl34_ = new_n_n367_ | new_n_n368_ | new_n_n369_;
  assign new_n_n1092_ = new_n_n475_ & new_ni3_;
  assign new_n_n1085_ = new_n_n520_ & new_n_n471_;
  assign new_n_n86_ = ~new_nw43_;
  assign new_n_n71_ = ~new_ni39_;
  assign new_n_n60_ = ~new_na33_;
  assign new_n_n53_ = ~new_nc31_;
  assign new_n_n42_ = ~new_nr28_;
  assign new_nh20_ = new_nl1_ & new_n_n337_ & new_n_n268_ & new_n_n361_;
  assign new_n_n1349_ = new_n_n356_ & new_nr1_ & new_np22_;
  assign new_na22_ = new_nf21_ | new_np22_;
  assign new_n_n1303_ = new_n_n363_ & new_n_n362_ & new_nt22_;
  assign new_n_n1295_ = new_n_n386_ & new_n_n243_;
  assign new_nw23_ = new_n_n1285_ | new_n_n1284_ | new_n_n1283_;
  assign new_na24_ = new_n_n1278_ | new_n_n1279_;
  assign new_ni24_ = new_nt23_ & new_nv1_;
  assign new_n_n1271_ = new_n_n212_ & new_n_n237_;
  assign new_n_n1244_ = new_n_n388_ & new_np25_;
  assign new_n_n1227_ = new_n_n241_ & new_n_n452_;
  assign new_n_n1223_ = new_nc2_ & new_nb2_;
  assign new_nu26_ = new_n_n1218_ | new_n_n1219_;
  assign new_n_n1213_ = new_n_n359_ & new_n_n253_;
  assign new_n_n1197_ = new_n_n257_ & new_n_n271_;
  assign new_na28_ = new_nm27_ & new_nk2_;
  assign new_n_n1186_ = new_nl2_ & new_n_n262_;
  assign new_nz28_ = new_n_n1170_ | new_n_n1171_;
  assign new_nf29_ = new_n_n1166_ | new_nh29_;
  assign new_n_n1162_ = new_n_n283_ & new_nt2_;
  assign new_n_n1157_ = new_n_n279_ & new_ne19_;
  assign new_nk30_ = new_n_n415_ | new_n_n365_ | new_n_n390_ | new_n_n340_;
  assign new_nx30_ = new_n_n1148_ | new_n_n1147_ | new_n_n1146_;
  assign new_n_n1143_ = new_n_n293_ & new_ne19_;
  assign new_n_n1137_ = new_n_n296_ & new_n_n324_;
  assign new_n_n1123_ = new_na3_ & new_n_n307_;
  assign new_ni33_ = new_nr20_ & new_n_n330_;
  assign new_ns33_ = new_n_n338_ | new_n_n445_;
  assign new_nb34_ = new_n_n357_ | new_n_n433_;
  assign new_nk34_ = new_n_n366_ | new_n_n451_;
  assign new_nf37_ = new_n_n1090_ | new_n_n1091_;
  assign new_n_n1086_ = new_nj50_ & new_n_n470_;
  assign new_n_n87_ = ~new_nj44_;
  assign new_n_n70_ = ~new_nu38_;
  assign new_n_n61_ = ~new_ng33_;
  assign new_n_n52_ = ~new_ny30_;
  assign new_n_n43_ = ~new_nv28_;
  assign new_ns5_ = ~new_ns35_;
  assign new_nf10_ = new_n_n111_ & new_n_n110_;
  assign new_nt10_ = new_n_n676_ & new_na53_;
  assign new_nm16_ = new_nu19_ & new_n_n136_;
  assign new_ne20_ = new_nw0_ & new_n_n356_;
  assign new_n_n1350_ = new_n_n356_ & new_nr1_ & new_nv20_;
  assign new_nm22_ = new_n_n268_ & new_n_n337_;
  assign new_n_n1305_ = new_n_n363_ & new_n_n362_ & new_n_n202_;
  assign new_n_n1296_ = new_ns1_ & new_nd21_;
  assign new_nu24_ = new_n_n1264_ | new_n_n1263_ | new_n_n1262_;
  assign new_nx24_ = new_n_n243_ & new_n_n221_;
  assign new_n_n1249_ = new_n_n225_ & new_nk20_;
  assign new_n_n1245_ = new_ny1_ & new_n_n229_;
  assign new_n_n1226_ = new_n_n242_ & new_n_n452_;
  assign new_n_n1221_ = new_nd2_ & new_nh26_;
  assign new_n_n1216_ = new_n_n250_ & new_n_n386_;
  assign new_nj27_ = new_nf27_ & new_ni2_;
  assign new_n_n1201_ = new_ni2_ & new_n_n256_;
  assign new_n_n1193_ = new_n_n259_ & new_n_n412_;
  assign new_nf28_ = new_n_n1185_ | new_n_n1186_;
  assign new_n_n1171_ = new_nq2_ & new_nr20_;
  assign new_n_n1165_ = new_n_n273_ & new_n_n414_;
  assign new_n_n1159_ = new_nr2_ & new_nt29_;
  assign new_nz29_ = new_n_n1151_ | new_n_n1152_;
  assign new_na30_ = new_n_n285_ | new_n_n284_;
  assign new_ns30_ = new_nv2_ & new_nq29_;
  assign new_n_n1144_ = new_n_n340_ & new_n_n290_;
  assign new_n_n1138_ = new_n_n297_ & new_ne19_;
  assign new_n_n1122_ = new_n_n450_ & new_nb32_;
  assign new_nh32_ = new_nr20_ & new_n_n314_;
  assign new_nv32_ = new_n_n1112_ | new_n_n1113_;
  assign new_na33_ = new_n_n322_ | new_n_n328_;
  assign new_nj34_ = new_n_n365_ | new_n_n449_;
  assign new_ni36_ = new_n_n1100_ | new_n_n1101_;
  assign new_nr36_ = new_n_n1094_ | new_n_n1095_;
  assign new_nn47_ = new_nr4_ & new_nt4_ & new_ny50_ & new_ns4_;
  assign new_nw47_ = new_n_n898_ | new_n_n899_;
  assign new_n_n830_ = new_n_n711_ & new_nw53_ & new_nx53_;
  assign new_n_n820_ = new_n_n711_ & new_n_n710_ & new_n_n678_;
  assign new_n_n797_ = ~new_nl0_;
  assign new_n_n88_ = ~new_nl44_;
  assign new_n_n33_ = ~new_no27_;
  assign new_n_n22_ = ~new_nr24_;
  assign new_n_n11_ = ~new_np18_;
  assign new_n_n0_ = ~new_nr16_;
  assign new_nt6_ = new_n_n268_ & new_nv21_;
  assign new_ne10_ = new_n_n111_ & new_n_n109_;
  assign new_nu10_ = new_n_n676_ & new_nc53_;
  assign new_nj16_ = new_n_n432_ | new_n_n381_ | new_n_n406_ | new_n_n356_;
  assign new_nf20_ = new_ng19_ & new_nv0_;
  assign new_n_n1351_ = new_np22_ & new_nh22_;
  assign new_n_n1323_ = new_n_n362_ & new_n_n363_;
  assign new_n_n1304_ = new_n_n362_ & new_nt22_ & new_n_n202_;
  assign new_ng23_ = new_n_n1295_ | new_n_n1296_;
  assign new_n_n1264_ = new_n_n218_ & new_nv19_;
  assign new_n_n1257_ = new_n_n220_ & new_nk20_;
  assign new_nc25_ = new_n_n243_ & new_n_n226_;
  assign new_nn25_ = new_n_n1244_ | new_n_n1245_;
  assign new_n_n1225_ = new_n_n242_ & new_nk20_;
  assign new_nm26_ = new_n_n1220_ | new_n_n1221_;
  assign new_n_n1209_ = new_ng2_ & new_nj26_;
  assign new_nm27_ = new_n_n1207_ | new_nl_;
  assign new_nq27_ = new_n_n1200_ | new_n_n1201_;
  assign new_n_n1192_ = new_n_n259_ & new_n_n271_;
  assign new_n_n1187_ = new_n_n261_ & new_n_n271_;
  assign new_n_n1170_ = new_n_n364_ & new_n_n285_;
  assign new_ng29_ = new_n_n1164_ | new_n_n1165_;
  assign new_n_n1158_ = new_n_n389_ & new_n_n276_;
  assign new_nx29_ = new_nr20_ & new_n_n281_;
  assign new_nb30_ = new_n_n1149_ | new_n_n1150_;
  assign new_nr30_ = new_nq29_ & new_nw2_;
  assign new_nz30_ = new_nr20_ & new_n_n291_;
  assign new_nf31_ = new_n_n1138_ | new_n_n1137_ | new_n_n1136_;
  assign new_nz31_ = new_n_n308_ | new_n_n328_;
  assign new_nf32_ = new_n_n313_ | new_n_n328_;
  assign new_n_n1113_ = new_nc3_ & new_nw32_;
  assign new_n_n1107_ = new_n_n416_ & new_nc33_;
  assign new_nz33_ = new_n_n355_ & new_n_n354_ & new_n_n353_;
  assign new_n_n1101_ = new_nf3_ & new_nc52_;
  assign new_n_n1096_ = new_nf3_ & new_ng3_;
  assign new_no47_ = new_n_n904_ | new_ni47_;
  assign new_n_n900_ = new_n_n600_ & new_n_n754_;
  assign new_n_n829_ = new_n_n710_ & new_n_n677_ & new_nx53_;
  assign new_n_n821_ = new_n_n711_ & new_n_n677_ & new_nx53_;
  assign new_n_n807_ = ~new_nv56_;
  assign new_n_n89_ = ~new_nw44_;
  assign new_n_n32_ = ~new_nd27_;
  assign new_n_n23_ = ~new_nw24_;
  assign new_n_n10_ = ~new_nm18_;
  assign new_n_n1_ = ~new_nu16_;
  assign new_ne7_ = new_nb_ | new_n_n24_;
  assign new_nj10_ = new_ne5_ | new_n_n114_;
  assign new_nr10_ = new_n_n121_ & new_n_n122_;
  assign new_n_n1380_ = new_n_n172_ & new_n_n362_;
  assign new_n_n1355_ = new_n_n164_ & new_nj1_;
  assign new_n_n1352_ = new_nh22_ & new_nv20_;
  assign new_n_n1315_ = new_n_n363_ & new_nt22_ & new_nu22_;
  assign new_n_n1263_ = new_n_n217_ & new_n_n237_;
  assign new_n_n1256_ = new_n_n223_ & new_nv19_;
  assign new_n_n1251_ = new_n_n241_ & new_n_n366_;
  assign new_n_n1246_ = new_n_n227_ & new_n_n228_;
  assign new_na26_ = new_n_n243_ & new_n_n244_;
  assign new_nv26_ = new_n_n1217_ | new_n_n1216_ | new_n_n1215_;
  assign new_nd27_ = new_n_n1208_ | new_n_n1209_;
  assign new_n_n1207_ = new_nj2_ & new_ni2_ & new_nf27_;
  assign new_nr27_ = new_n_n1199_ | new_n_n1198_ | new_n_n1197_;
  assign new_nu27_ = new_n_n1194_ | new_n_n1193_ | new_n_n1192_;
  assign new_n_n1188_ = new_n_n261_ & new_n_n444_;
  assign new_nc29_ = new_n_n1169_ | new_nh29_;
  assign new_nh29_ = new_n_n274_ & new_n_n275_;
  assign new_n_n1160_ = new_n_n324_ & new_n_n364_;
  assign new_n_n1153_ = new_n_n414_ & new_n_n280_;
  assign new_n_n1150_ = new_nt2_ & new_na30_;
  assign new_nu30_ = new_nx2_ & new_nw2_ & new_nq29_;
  assign new_ny30_ = new_n_n1144_ | new_n_n1145_;
  assign new_nd31_ = new_nr20_ & new_n_n295_;
  assign new_nb32_ = new_nr20_ & new_n_n309_;
  assign new_np32_ = new_ne3_ | new_nc3_ | new_nd3_ | new_nb3_;
  assign new_n_n1115_ = new_np31_ & new_n_n324_;
  assign new_n_n1108_ = new_nd3_ & new_n_n321_;
  assign new_np33_ = new_no28_ | new_n_n439_;
  assign new_nn35_ = new_n_n415_ | new_n_n449_;
  assign new_ny35_ = new_n_n442_ | new_n_n441_;
  assign new_ng44_ = new_nd4_ & new_ne4_;
  assign new_nj47_ = new_ny50_ & new_n_n605_;
  assign new_n_n901_ = new_nl47_ & new_nt4_;
  assign new_np53_ = new_nm53_ | new_n_n670_;
  assign new_n_n837_ = new_n_n710_ & new_n_n686_;
  assign new_na57_ = new_n_n796_ | new_n_n795_;
  assign new_n_n31_ = ~new_nz26_;
  assign new_n_n20_ = ~new_nw23_;
  assign new_n_n13_ = ~new_nb20_;
  assign new_n_n2_ = ~new_nw16_;
  assign new_no7_ = new_nb_ | new_n_n33_;
  assign new_ng10_ = new_n_n111_ & new_n_n112_;
  assign new_ns10_ = new_n_n676_ & new_nk53_;
  assign new_n_n1381_ = new_n_n172_ & new_nh22_;
  assign new_nc20_ = new_no19_ & new_n_n181_;
  assign new_nn20_ = new_n_n1349_ | new_n_n1351_ | new_n_n1350_ | new_n_n1352_;
  assign new_n_n1306_ = new_n_n363_ & new_n_n201_ & new_nu22_;
  assign new_n_n1262_ = new_n_n217_ & new_n_n218_;
  assign new_nz24_ = new_n_n1256_ | new_n_n1255_ | new_n_n1254_;
  assign new_n_n1250_ = new_n_n225_ & new_n_n366_;
  assign new_n_n1247_ = new_n_n227_ & new_n_n237_;
  assign new_n_n1220_ = new_n_n408_ & new_n_n246_;
  assign new_n_n1217_ = new_nq19_ & new_n_n386_;
  assign new_n_n1210_ = new_n_n251_ & new_n_n271_;
  assign new_nn27_ = new_n_n1205_ | new_n_n1206_;
  assign new_n_n1200_ = new_n_n409_ & new_nf27_;
  assign new_n_n1194_ = new_nq19_ & new_n_n412_;
  assign new_n_n1189_ = new_nq19_ & new_n_n444_;
  assign new_n_n1169_ = new_n_n364_ & new_n_n389_;
  assign new_n_n1164_ = new_n_n273_ & new_n_n278_;
  assign new_ns29_ = new_n_n1158_ | new_n_n1159_;
  assign new_n_n1154_ = new_ns2_ & new_nx29_;
  assign new_n_n1149_ = new_n_n448_ & new_n_n286_;
  assign new_nt30_ = new_nn29_ & new_n_n340_ & new_n_n365_;
  assign new_n_n1145_ = new_nw2_ & new_nz30_;
  assign new_n_n1139_ = new_n_n365_ & new_n_n294_;
  assign new_nd32_ = new_n_n1121_ | new_n_n1120_ | new_n_n1119_;
  assign new_nl32_ = new_n_n390_ | new_nz2_ | new_na3_;
  assign new_n_n1114_ = new_np31_ & new_nn31_;
  assign new_nz32_ = new_n_n1107_ | new_n_n1108_;
  assign new_nf33_ = new_n_n1102_ | new_n_n1103_;
  assign new_no35_ = new_n_n416_ | new_n_n451_;
  assign new_nx35_ = new_n_n440_ | new_n_n439_;
  assign new_nr44_ = new_n_n577_ | new_n_n784_;
  assign new_nl47_ = new_nr4_ & new_ns4_ & new_ny50_;
  assign new_nt47_ = new_n_n900_ | new_n_n901_;
  assign new_nq53_ = new_nm5_ & new_nl5_;
  assign new_n_n838_ = new_n_n710_ & new_n_n711_;
  assign new_nq56_ = new_n_n775_ | new_n_n773_ | new_n_n774_ | new_n_n772_;
  assign new_n_n30_ = ~new_nv26_;
  assign new_n_n21_ = ~new_nb24_;
  assign new_n_n12_ = ~new_nq18_;
  assign new_n_n3_ = ~new_nz16_;
  assign new_n_n1389_ = new_nb16_ & new_np2_;
  assign new_nu16_ = new_n_n1377_ | new_n_n1378_;
  assign new_ne17_ = new_nu19_ & new_nc1_;
  assign new_nr17_ = new_n_n1367_ | new_n_n1368_;
  assign new_nc18_ = new_n_n1361_ | new_n_n1362_;
  assign new_n_n1344_ = new_n_n362_ & new_n_n168_ & new_n_n338_;
  assign new_nd21_ = new_n_n176_ & new_n_n177_;
  assign new_n_n1334_ = new_n_n197_ & new_np21_;
  assign new_n_n1327_ = new_nh22_ & new_n_n361_ & new_n_n197_;
  assign new_ni22_ = new_nr18_ | new_n_n194_;
  assign new_nu22_ = new_n_n199_ & new_n_n200_;
  assign new_n_n1317_ = new_n_n338_ & new_n_n362_ & new_n_n201_;
  assign new_n_n1307_ = new_n_n338_ & new_nt22_ & new_nu22_;
  assign new_n_n1278_ = new_n_n442_ & new_nc24_;
  assign new_n_n1274_ = new_n_n444_ & new_n_n387_ & new_nr23_ & new_n_n412_;
  assign new_n_n1267_ = new_n_n241_ & new_n_n415_;
  assign new_nw24_ = new_n_n1259_ | new_n_n1258_ | new_n_n1257_;
  assign new_n_n1252_ = new_n_n444_ & new_nc25_;
  assign new_n_n1248_ = new_n_n228_ & new_nv19_;
  assign new_n_n1238_ = new_n_n232_ & new_n_n233_;
  assign new_n_n1204_ = new_nq19_ & new_n_n442_;
  assign new_n_n1196_ = new_nj2_ & new_n_n258_;
  assign new_nd28_ = new_n_n1189_ | new_n_n1188_ | new_n_n1187_;
  assign new_nj28_ = new_n_n1179_ | new_n_n1178_ | new_n_n1177_;
  assign new_n_n1176_ = new_no2_ & new_n_n269_;
  assign new_no31_ = new_n_n1132_ | new_nj_;
  assign new_nv31_ = new_nr20_ & new_n_n304_;
  assign new_nt34_ = new_n_n385_ | new_n_n439_;
  assign new_ne35_ = new_n_n406_ | new_n_n431_;
  assign new_nz44_ = new_n_n948_ | new_n_n949_;
  assign new_nf48_ = new_n_n605_ & new_nv4_ & new_ny50_;
  assign new_n_n892_ = new_n_n608_ & new_n_n730_;
  assign new_n_n886_ = new_n_n611_ & new_no49_;
  assign new_nr49_ = new_n_n620_ | new_n_n628_;
  assign new_nw52_ = new_n_n846_ | new_n_n847_;
  assign new_nc53_ = new_n_n661_ | new_n_n660_;
  assign new_ng56_ = new_n_n757_ | new_n_n785_;
  assign new_n_n59_ = ~new_nv32_;
  assign new_n_n48_ = ~new_nw29_;
  assign new_n_n37_ = ~new_ng28_;
  assign new_n_n26_ = ~new_nt25_;
  assign new_n_n15_ = ~new_nz22_;
  assign new_n_n4_ = ~new_nm17_;
  assign new_nc8_ = new_n_n51_ & new_nt20_;
  assign new_n_n1378_ = new_nl16_ & new_nw0_;
  assign new_nd17_ = new_n_n135_ & new_n_n136_;
  assign new_n_n1368_ = new_nl17_ & new_nb1_;
  assign new_nb18_ = new_nb_ | new_n_n159_;
  assign new_n_n1343_ = new_n_n169_ & new_n_n168_ & new_n_n338_;
  assign new_nc21_ = new_n_n175_ & new_nv6_;
  assign new_n_n1333_ = new_n_n197_ & new_n_n339_;
  assign new_n_n1328_ = new_np21_ & new_n_n337_ & new_n_n197_;
  assign new_nj22_ = new_np21_ | new_nr18_ | new_n_n339_;
  assign new_nt22_ = new_n_n197_ & new_n_n198_;
  assign new_n_n1316_ = new_n_n363_ & new_n_n362_ & new_nu22_;
  assign new_n_n1308_ = new_n_n363_ & new_n_n338_ & new_nu22_;
  assign new_nb24_ = new_n_n1277_ | new_n_n1276_ | new_n_n1275_;
  assign new_nm24_ = new_n_n1274_ | new_nk_;
  assign new_n_n1266_ = new_n_n215_ & new_n_n415_;
  assign new_n_n1260_ = new_n_n412_ & new_nx24_;
  assign new_nb25_ = new_n_n1251_ | new_n_n1250_ | new_n_n1249_;
  assign new_nm25_ = new_n_n1248_ | new_n_n1247_ | new_n_n1246_;
  assign new_n_n1232_ = new_n_n239_ & new_nv19_;
  assign new_n_n1208_ = new_n_n436_ & new_n_n252_;
  assign new_n_n1195_ = new_n_n438_ & new_nj27_;
  assign new_n_n1190_ = new_n_n360_ & new_nm27_;
  assign new_n_n1179_ = new_nq19_ & new_n_n413_;
  assign new_nu28_ = new_n_n1175_ | new_n_n1176_;
  assign new_n_n1132_ = new_ns30_ & new_na3_;
  assign new_nt31_ = new_n_n303_ | new_n_n328_;
  assign new_nu34_ = new_n_n386_ | new_n_n441_;
  assign new_nd35_ = new_n_n405_ & new_n_n404_ & new_n_n403_;
  assign new_ng45_ = new_nj4_ & new_nh4_ & new_n_n578_;
  assign new_ng48_ = new_n_n605_ & new_n_n604_ & new_ny50_;
  assign new_n_n893_ = new_ni48_ & new_nx4_;
  assign new_nb49_ = new_n_n884_ | new_n_n885_;
  assign new_np49_ = new_n_n618_ & new_n_n619_;
  assign new_n_n847_ = new_nm53_ & new_n_n656_ & new_n_n674_;
  assign new_na53_ = new_n_n659_ | new_n_n658_;
  assign new_nw55_ = new_n_n737_ | new_n_n795_;
  assign new_n_n58_ = ~new_nf32_;
  assign new_n_n49_ = ~new_nc30_;
  assign new_n_n36_ = ~new_nd28_;
  assign new_n_n27_ = ~new_ny25_;
  assign new_n_n14_ = ~new_nc20_;
  assign new_n_n5_ = ~new_no17_;
  assign new_nm8_ = new_ne52_ & new_n_n62_;
  assign new_n_n1377_ = new_n_n130_ & new_n_n381_;
  assign new_ni17_ = new_n_n136_ & new_nz0_ & new_nu19_;
  assign new_n_n1370_ = new_ni17_ & new_na1_;
  assign new_n_n1363_ = new_n_n141_ & new_nd1_;
  assign new_n_n1342_ = new_n_n362_ & new_n_n363_ & new_n_n338_;
  assign new_nf21_ = new_n_n1339_ | new_n_n1338_ | new_n_n1337_;
  assign new_n_n1336_ = new_n_n197_ & new_nh22_;
  assign new_n_n1329_ = new_n_n182_ & new_n_n337_ & new_n_n197_;
  assign new_nk22_ = new_nh22_ | new_n_n195_;
  assign new_n_n1324_ = new_n_n338_ & new_n_n363_;
  assign new_nc23_ = new_n_n1316_ | new_n_n1315_ | new_n_n1318_ | new_n_n1317_ | new_n_n1314_ | new_n_n1313_ | new_n_n1311_ | new_n_n1312_;
  assign new_n_n1309_ = new_n_n363_ & new_n_n362_ & new_n_n201_;
  assign new_n_n1291_ = new_n_n442_ & new_n_n411_ & new_n_n386_;
  assign new_n_n1284_ = new_n_n205_ & new_n_n365_;
  assign new_n_n1265_ = new_n_n215_ & new_nk20_;
  assign new_n_n1258_ = new_n_n220_ & new_n_n450_;
  assign new_na25_ = new_n_n1252_ | new_n_n1253_;
  assign new_nl25_ = new_nz1_ & new_ny1_ & new_no24_;
  assign new_n_n1240_ = new_n_n233_ & new_nv19_;
  assign new_nw25_ = new_n_n1232_ | new_n_n1231_ | new_n_n1230_;
  assign new_nf27_ = new_nh2_ & new_nf2_ & new_n_n253_;
  assign new_n_n1202_ = new_n_n255_ & new_n_n271_;
  assign new_n_n1191_ = new_nk2_ & new_n_n260_;
  assign new_n_n1181_ = new_nm2_ & new_n_n264_;
  assign new_nt28_ = new_n_n268_ & new_nq19_;
  assign new_n_n1133_ = new_nq30_ & new_n_n450_;
  assign new_n_n1127_ = new_n_n415_ & new_nv31_;
  assign new_n_n938_ = new_nv50_ & new_n_n790_;
  assign new_ni48_ = new_n_n605_ & new_nw4_ & new_ny50_ & new_nv4_;
  assign new_n_n891_ = new_ng48_ & new_ny4_;
  assign new_nz48_ = new_n_n886_ | new_n_n887_;
  assign new_no49_ = new_nb5_ | new_n_n617_;
  assign new_n_n856_ = new_n_n647_ & new_n_n648_;
  assign new_n_n853_ = new_n_n655_ & new_n_n782_ & new_ns48_;
  assign new_nm55_ = new_n_n725_ | new_n_n723_ | new_n_n724_ | new_n_n722_;
  assign new_n_n79_ = ~new_nu41_;
  assign new_n_n68_ = ~new_nm38_;
  assign new_n_n35_ = ~new_nu27_;
  assign new_n_n24_ = ~new_nb25_;
  assign new_n_n17_ = ~new_nd23_;
  assign new_n_n6_ = ~new_nr17_;
  assign new_nt8_ = new_ne52_ & new_n_n69_;
  assign new_nw16_ = new_n_n1375_ | new_n_n1376_;
  assign new_nf17_ = new_n_n335_ | new_n_n357_ | new_n_n382_;
  assign new_n_n1369_ = new_n_n138_ & new_n_n357_;
  assign new_n_n1364_ = new_nb17_ & new_n_n434_;
  assign new_n_n1341_ = new_n_n169_ & new_n_n363_ & new_n_n338_;
  assign new_ne21_ = new_n_n334_ & new_n_n337_ & new_n_n268_ & new_nm1_;
  assign new_n_n1335_ = new_n_n197_ & new_nr18_;
  assign new_n_n1330_ = new_nh22_ & new_n_n337_ & new_n_n197_;
  assign new_nl22_ = new_nm1_ & new_nl1_;
  assign new_nv22_ = new_n_n1324_ | new_n_n1323_ | new_n_n1322_;
  assign new_n_n1318_ = new_n_n363_ & new_n_n338_ & new_nt22_;
  assign new_n_n1310_ = new_n_n338_ & new_n_n362_ & new_nt22_;
  assign new_nt23_ = new_n_n1290_ | new_nk_;
  assign new_n_n1285_ = new_n_n241_ & new_n_n365_;
  assign new_ns24_ = new_n_n243_ & new_n_n216_;
  assign new_n_n1259_ = new_n_n241_ & new_n_n450_;
  assign new_n_n1253_ = new_nx1_ & new_n_n224_;
  assign new_nj25_ = new_nm24_ & new_n_n388_ & new_n_n413_;
  assign new_n_n1239_ = new_n_n232_ & new_n_n237_;
  assign new_nu25_ = new_n_n243_ & new_n_n236_;
  assign new_nh27_ = new_n_n253_ & new_nf2_;
  assign new_n_n1203_ = new_n_n255_ & new_n_n442_;
  assign new_nt27_ = new_n_n1195_ | new_n_n1196_;
  assign new_n_n1180_ = new_n_n410_ & new_nx27_;
  assign new_ns28_ = new_nx27_ & new_nm2_;
  assign new_nn31_ = new_nb3_ | new_n_n311_;
  assign new_n_n1128_ = new_nz2_ & new_n_n302_;
  assign new_n_n931_ = new_nl4_ & new_n_n583_;
  assign new_nj48_ = new_n_n896_ | new_n_n897_;
  assign new_nq48_ = new_n_n890_ | new_n_n891_;
  assign new_n_n887_ = new_n_n611_ & new_n_n623_;
  assign new_nn49_ = new_n_n624_ | new_n_n616_;
  assign new_nc52_ = new_nd0_ | new_n_n649_;
  assign new_n_n854_ = new_n_n655_ & new_n_n782_ & new_n_n710_;
  assign new_nc55_ = new_n_n707_ | new_n_n785_;
  assign new_n_n78_ = ~new_ne41_;
  assign new_n_n69_ = ~new_nq38_;
  assign new_n_n34_ = ~new_nr27_;
  assign new_n_n25_ = ~new_no25_;
  assign new_n_n16_ = ~new_nc23_;
  assign new_n_n7_ = ~new_nt17_;
  assign new_nd9_ = new_n_n676_ & new_n_n80_;
  assign new_nl18_ = new_n_n146_ | new_n_n145_ | new_nu18_;
  assign new_n_n1357_ = new_n_n156_ & new_nr18_;
  assign new_nz19_ = new_nj1_ | new_no1_;
  assign new_nr20_ = new_nf_ | new_n_n170_;
  assign new_n_n1338_ = new_n_n178_ & new_n_n434_ & new_nv17_;
  assign new_nr21_ = new_n_n1331_ | new_n_n1332_;
  assign new_nx21_ = new_n_n186_ | new_n_n185_;
  assign new_nc22_ = new_n_n188_ | new_n_n187_;
  assign new_nq22_ = new_n_n361_ & new_n_n334_;
  assign new_n_n1320_ = new_nr1_ & new_nv22_ & new_n_n268_;
  assign new_n_n1311_ = new_n_n363_ & new_n_n338_ & new_n_n362_;
  assign new_n_n1298_ = new_n_n363_ & new_n_n338_ & new_n_n202_;
  assign new_nr23_ = new_n_n1291_ | new_nk_;
  assign new_n_n1290_ = new_nu1_ & new_nt1_ & new_ns1_;
  assign new_nx23_ = new_n_n243_ & new_n_n206_;
  assign new_n_n1275_ = new_n_n210_ & new_nk20_;
  assign new_n_n1272_ = new_n_n213_ & new_nv19_;
  assign new_n_n1255_ = new_n_n222_ & new_n_n237_;
  assign new_ni25_ = new_no24_ & new_ny1_;
  assign new_np25_ = new_n_n243_ & new_n_n231_;
  assign new_n_n1233_ = new_n_n235_ & new_nk20_;
  assign new_nf26_ = new_nl_ | new_n_n338_;
  assign new_nr26_ = new_n_n252_ | new_n_n436_;
  assign new_n_n1214_ = new_nf2_ & new_no26_;
  assign new_n_n1182_ = new_n_n263_ & new_n_n271_;
  assign new_nr28_ = new_n_n440_ | new_n_n410_ | new_n_n385_;
  assign new_ns31_ = new_n_n1127_ | new_n_n1128_;
  assign new_n_n925_ = new_n_n708_ & new_nn45_;
  assign new_nz49_ = new_n_n630_ & new_n_n628_;
  assign new_nl50_ = new_nn50_ & new_n_n729_ & new_n_n782_;
  assign new_n_n875_ = new_np46_ & new_n_n637_;
  assign new_np51_ = new_n_n868_ | new_n_n870_ | new_n_n869_ | new_n_n871_;
  assign new_n_n871_ = new_nf52_ & new_n_n640_;
  assign new_n_n861_ = new_n_n710_ & new_n_n643_ & new_n_n642_;
  assign new_ns54_ = new_n_n687_ | new_n_n795_;
  assign new_n_n80_ = ~new_nz41_;
  assign new_n_n77_ = ~new_nx40_;
  assign new_n_n66_ = ~new_nt37_;
  assign new_n_n55_ = ~new_nt31_;
  assign new_n_n44_ = ~new_nb16_;
  assign new_n_n19_ = ~new_ni23_;
  assign new_n_n8_ = ~new_ns16_;
  assign new_nn9_ = new_nz_ | new_n_n89_;
  assign new_nm18_ = new_n_n154_ | new_n_n144_;
  assign new_n_n1358_ = new_nu18_ & new_n_n182_;
  assign new_nb20_ = new_nb_ | new_n_n1356_ | new_n_n1355_;
  assign new_nt20_ = new_n_n194_ & new_n_n268_;
  assign new_n_n1339_ = new_n_n178_ & new_n_n434_ & new_n_n362_;
  assign new_n_n1332_ = new_nh22_ & new_n_n181_ & new_n_n199_;
  assign new_nv21_ = new_n_n184_ | new_n_n183_;
  assign new_nd22_ = new_n_n189_ & new_n_n194_ & new_n_n199_;
  assign new_np22_ = new_n_n268_ & new_nn22_;
  assign new_n_n1319_ = new_nq1_ & new_nv22_ & new_n_n268_;
  assign new_nd23_ = new_n_n1308_ | new_n_n1307_ | new_n_n1310_ | new_n_n1309_ | new_n_n1306_ | new_n_n1305_ | new_n_n1311_ | new_n_n1304_;
  assign new_n_n1297_ = new_n_n363_ & new_nt22_ & new_n_n202_;
  assign new_nq23_ = new_ns1_ & new_nt1_;
  assign new_nu23_ = new_n_n1288_ | new_n_n1289_;
  assign new_n_n1283_ = new_n_n205_ & new_nk20_;
  assign new_nc24_ = new_n_n243_ & new_n_n211_;
  assign new_np24_ = new_n_n1272_ | new_n_n1271_ | new_n_n1270_;
  assign new_n_n1254_ = new_n_n222_ & new_n_n223_;
  assign new_ng25_ = new_n_n388_ & new_nm24_;
  assign new_nr25_ = new_n_n1240_ | new_n_n1239_ | new_n_n1238_;
  assign new_n_n1234_ = new_n_n235_ & new_n_n416_;
  assign new_n_n1231_ = new_n_n238_ & new_n_n237_;
  assign new_ns26_ = new_n_n363_ & new_n_n247_;
  assign new_ny26_ = new_n_n1213_ | new_n_n1214_;
  assign new_ni28_ = new_n_n1180_ | new_n_n1181_;
  assign new_nq28_ = new_n_n360_ | new_n_n438_ | new_n_n409_;
  assign new_nl31_ = new_n_n1133_ | new_nj_;
  assign new_n_n918_ = new_nv50_ & new_n_n736_;
  assign new_na50_ = new_n_n881_ | new_n_n880_ | new_n_n879_;
  assign new_nj50_ = new_n_n631_ & new_n_n632_;
  assign new_n_n874_ = new_n_n638_ & new_nh5_;
  assign new_nm51_ = new_n_n645_ & new_nk5_;
  assign new_n_n870_ = new_nu53_ & new_n_n640_;
  assign new_n_n862_ = new_n_n711_ & new_n_n644_ & new_n_n642_;
  assign new_n_n812_ = new_n_n711_ & new_nw53_ & new_n_n678_;
  assign new_n_n81_ = ~new_np42_;
  assign new_n_n76_ = ~new_nr40_;
  assign new_n_n67_ = ~new_ny37_;
  assign new_n_n54_ = ~new_ng31_;
  assign new_n_n45_ = ~new_na_;
  assign new_n_n18_ = ~new_ne23_;
  assign new_n_n9_ = ~new_ny17_;
  assign new_nx9_ = new_nz_ | new_n_n102_;
  assign new_np18_ = new_nr18_ | new_n_n145_ | new_n_n146_;
  assign new_ng19_ = new_ni19_ & new_n_n381_ & new_n_n434_;
  assign new_nv19_ = new_n_n172_ & new_n_n161_;
  assign new_n_n1354_ = new_n_n181_ & new_n_n165_;
  assign new_nv20_ = new_n_n1340_ | new_n_n171_;
  assign new_nm21_ = new_ne3_ & new_nd3_ & new_nc3_;
  assign new_np21_ = new_n_n179_ & new_n_n180_;
  assign new_n_n1325_ = new_np21_ & new_n_n361_ & new_n_n197_;
  assign new_nf22_ = new_n_n190_ | new_nh20_ | new_n_n191_;
  assign new_ns22_ = new_n_n338_ | new_nh22_;
  assign new_nz22_ = new_n_n1321_ | new_n_n1320_ | new_n_n1319_;
  assign new_n_n1312_ = new_n_n338_ & new_nt22_ & new_n_n202_;
  assign new_n_n1300_ = new_n_n362_ & new_nt22_ & new_nu22_;
  assign new_no23_ = new_n_n411_ & new_n_n386_;
  assign new_n_n1289_ = new_nv19_ & new_ns1_;
  assign new_n_n1282_ = new_n_n208_ & new_nv19_;
  assign new_n_n1277_ = new_n_n241_ & new_n_n390_;
  assign new_n_n1273_ = new_nx1_ & new_nv1_ & new_nt23_ & new_nw1_;
  assign new_n_n1268_ = new_n_n387_ & new_ns24_;
  assign new_n_n1261_ = new_nw1_ & new_n_n219_;
  assign new_n_n1242_ = new_n_n230_ & new_n_n391_;
  assign new_n_n1235_ = new_n_n241_ & new_n_n416_;
  assign new_n_n1230_ = new_n_n238_ & new_n_n239_;
  assign new_nj26_ = new_n_n1224_ | new_n_n245_;
  assign new_n_n1215_ = new_n_n250_ & new_n_n271_;
  assign new_n_n1184_ = new_nq19_ & new_n_n388_;
  assign new_np28_ = new_n_n359_ | new_n_n384_;
  assign new_nr46_ = new_n_n707_ | new_n_n732_;
  assign new_n_n881_ = new_n_n676_ & new_n_n630_ & new_nx49_;
  assign new_np50_ = new_n_n780_ & new_n_n754_;
  assign new_nb51_ = new_ng5_ | new_no5_;
  assign new_n_n872_ = new_n_n656_ & new_nu53_;
  assign new_n_n82_ = ~new_nu42_;
  assign new_n_n75_ = ~new_nm40_;
  assign new_n_n64_ = ~new_nk37_;
  assign new_n_n57_ = ~new_nd30_;
  assign new_n_n46_ = ~new_nz28_;
  assign new_n_n39_ = ~new_nt28_;
  assign new_n_n28_ = ~new_nk26_;
  assign new_nq18_ = new_n_n155_ | new_n_n147_;
  assign new_ne19_ = new_n_n157_ & new_n_n158_;
  assign new_ny19_ = new_nk1_ | new_n_n162_;
  assign new_n_n1346_ = new_n_n362_ & new_n_n167_ & new_n_n363_;
  assign new_n_n1340_ = new_n_n172_ & new_n_n173_;
  assign new_n_n1337_ = new_n_n178_ & new_nr1_ & new_nv17_;
  assign new_nq21_ = new_n_n334_ & new_nn1_ & new_n_n268_ & new_n_n361_;
  assign new_n_n1326_ = new_n_n182_ & new_n_n361_ & new_n_n197_;
  assign new_nh22_ = new_n_n193_ | new_n_n192_;
  assign new_nr22_ = new_n_n363_ | new_nh22_;
  assign new_n_n1321_ = new_np1_ & new_nv22_ & new_n_n268_;
  assign new_n_n1313_ = new_n_n338_ & new_n_n362_ & new_n_n202_;
  assign new_n_n1299_ = new_n_n338_ & new_n_n201_ & new_nu22_;
  assign new_n_n1292_ = new_n_n203_ & new_nk20_;
  assign new_n_n1288_ = new_n_n237_ & new_n_n386_;
  assign new_nz23_ = new_n_n1282_ | new_n_n1281_ | new_n_n1280_;
  assign new_n_n1276_ = new_n_n210_ & new_n_n390_;
  assign new_no24_ = new_n_n1273_ | new_nk_;
  assign new_nr24_ = new_n_n1267_ | new_n_n1266_ | new_n_n1265_;
  assign new_nv24_ = new_n_n1260_ | new_n_n1261_;
  assign new_n_n1241_ = new_n_n230_ & new_nk20_;
  assign new_nt25_ = new_n_n1235_ | new_n_n1234_ | new_n_n1233_;
  assign new_nx25_ = new_n_n1228_ | new_n_n1229_;
  assign new_nh26_ = new_nb2_ & new_nc2_;
  assign new_no26_ = new_n_n266_ | new_n_n336_;
  assign new_n_n1183_ = new_n_n263_ & new_n_n388_;
  assign new_no28_ = new_n_n266_ | new_n_n336_ | new_n_n267_;
  assign new_n_n908_ = new_nv50_ & new_n_n794_;
  assign new_n_n880_ = new_n_n676_ & new_n_n630_ & new_n_n627_;
  assign new_nn50_ = new_nr50_ & new_n_n730_ & new_n_n755_ & new_n_n705_;
  assign new_nd51_ = new_nz_ | new_n_n875_ | new_n_n874_;
  assign new_n_n873_ = new_n_n656_ & new_n_n639_;
  assign new_n_n83_ = ~new_nz42_;
  assign new_n_n74_ = ~new_nu39_;
  assign new_n_n65_ = ~new_nq37_;
  assign new_n_n56_ = ~new_nz31_;
  assign new_n_n47_ = ~new_ns29_;
  assign new_n_n38_ = ~new_nj28_;
  assign new_n_n29_ = ~new_nm26_;
endmodule


