// Benchmark "top" written by ABC on Fri Mar 31 12:09:22 2023

module top ( 
    pdel1, pratr, pbull1, pbull0, pwatch, povacc, pverr_n, porwd_n,
    pvlenesr, pmmerr, paccrpy, pvacc, pcat4, pvst1, pcapsd, pcat3, pcat2,
    pcat1, plsd, pvst0, pcat0, pibt2, pkbg_n, pmarssr, pend, pvsumesr,
    pbull5, ppluto4, pstar2, pbull4, ppluto5, ppy, pstar3, pbull3,
    pcomppar, pibt1, pstar0, pbull2, pibt0, pstar1, ppluto0, pfbi, powl_n,
    ppluto1, piclr, ppluto2, pbull6, pcat5, ppluto3,
    pbull2_p, pend_p, pbull3_p, porwd_f, pbull4_p, ppluto3_p, pwatch_p,
    pbull5_p, pbull6_p, ppluto5_p, ppy_p, ppluto4_p, plsd_p, pvlenesr_p,
    pfbi_p, pstar1_p, pvsumesr_p, paccrpy_p, pkbg_f, pmarssr_p, pstar0_p,
    pstar3_p, pdel1_p, pstar2_p, pvst0_p, pcomppar_p, powl_f, psdo,
    pvst1_p, ppluto1_p, pratr_p, ppluto0_p, povacc_p, ppluto2_p, pbull0_p,
    pverr_f, pbull1_p  );
  input  pdel1, pratr, pbull1, pbull0, pwatch, povacc, pverr_n, porwd_n,
    pvlenesr, pmmerr, paccrpy, pvacc, pcat4, pvst1, pcapsd, pcat3, pcat2,
    pcat1, plsd, pvst0, pcat0, pibt2, pkbg_n, pmarssr, pend, pvsumesr,
    pbull5, ppluto4, pstar2, pbull4, ppluto5, ppy, pstar3, pbull3,
    pcomppar, pibt1, pstar0, pbull2, pibt0, pstar1, ppluto0, pfbi, powl_n,
    ppluto1, piclr, ppluto2, pbull6, pcat5, ppluto3;
  output pbull2_p, pend_p, pbull3_p, porwd_f, pbull4_p, ppluto3_p, pwatch_p,
    pbull5_p, pbull6_p, ppluto5_p, ppy_p, ppluto4_p, plsd_p, pvlenesr_p,
    pfbi_p, pstar1_p, pvsumesr_p, paccrpy_p, pkbg_f, pmarssr_p, pstar0_p,
    pstar3_p, pdel1_p, pstar2_p, pvst0_p, pcomppar_p, powl_f, psdo,
    pvst1_p, ppluto1_p, pratr_p, ppluto0_p, povacc_p, ppluto2_p, pbull0_p,
    pverr_f, pbull1_p;
  wire new_ndel1_, new_nratr_, new_nbull1_, new_nbull0_, new_nwatch_,
    new_novacc_, new_nverr_n_, new_norwd_n_, new_nvlenesr_, new_nmmerr_,
    new_naccrpy_, new_nvacc_, new_ncat4_, new_nvst1_, new_ncapsd_,
    new_ncat3_, new_ncat2_, new_ncat1_, new_nlsd_, new_nvst0_, new_ncat0_,
    new_nibt2_, new_nkbg_n_, new_nmarssr_, new_nend_, new_nvsumesr_,
    new_nbull5_, new_npluto4_, new_nstar2_, new_nbull4_, new_npluto5_,
    new_npy_, new_nstar3_, new_nbull3_, new_ncomppar_, new_nibt1_,
    new_nstar0_, new_nbull2_, new_nibt0_, new_nstar1_, new_npluto0_,
    new_nfbi_, new_nowl_n_, new_npluto1_, new_niclr_, new_npluto2_,
    new_nbull6_, new_ncat5_, new_npluto3_, new_naccrpy_p_, new_n_n119_,
    new_n_n111_, new_nvst1_p_, new_nstar2_p_, new_n_n87_, new_nbull4_p_,
    new_n_n147_, new_n_n118_, new_nkbg_f_, new_n_n103_, new_n_n96_,
    new_n_n86_, new_n_n80_, new_n_n148_, new_npluto3_p_, new_n_n125_,
    new_n_n102_, new_n_n94_, new_n_n88_, new_n_n81_, new_n_n149_,
    new_n_n131_, new_nowl_f_, new_nstar0_p_, new_n_n95_, new_nbull0_p_,
    new_nbull3_p_, new_n_n144_, new_npluto0_p_, new_n_n101_, new_n_n92_,
    new_n_n84_, new_nbull5_p_, new_n_n9_, new_n_n145_, new_n_n143_,
    new_n_n138_, new_n_n100_, new_n_n93_, new_nbull2_p_, new_n_n77_,
    new_nverr_f_, new_nstar1_p_, new_n_n91_, new_nbull1_p_, new_n_n78_,
    new_n_n146_, new_n_n99_, new_nstar3_p_, new_n_n85_, new_n_n79_,
    new_nmarssr_p_, new_n_n135_, new_npluto5_p_, new_n_n121_, new_n_n112_,
    new_nvst0_p_, new_n_n5_, new_n_n141_, new_npluto1_p_, new_n_n127_,
    new_nend_p_, new_novacc_p_, new_n_n106_, new_n_n6_, new_nratr_p_,
    new_n_n136_, new_n_n126_, new_n_n120_, new_n_n113_, new_n_n107_,
    new_n_n7_, new_n_n142_, new_n_n137_, new_norwd_f_, new_nfbi_p_,
    new_nwatch_p_, new_n_n108_, new_n_n8_, new_n_n150_, new_nvsumesr_p_,
    new_n_n132_, new_n_n130_, new_npy_p_, new_n_n115_, new_ncomppar_p_,
    new_n_n90_, new_n_n82_, new_n_n1_, new_nlsd_p_, new_n_n139_,
    new_n_n133_, new_npluto4_p_, new_n_n124_, new_n_n114_, new_ndel1_p_,
    new_n_n89_, new_n_n83_, new_n_n2_, new_nvlenesr_p_, new_npluto2_p_,
    new_n_n129_, new_n_n122_, new_n_n117_, new_n_n109_, new_n_n105_,
    new_n_n97_, new_n_n3_, new_n_n140_, new_n_n134_, new_n_n128_,
    new_n_n123_, new_n_n116_, new_n_n110_, new_n_n104_, new_n_n98_,
    new_n_n4_, new_n_n72_, new_n_n64_, new_n__1015_m__, new_n_n51_,
    new_n_n48_, new_nbull6_p_, new_n__219_m__, new_nc29g7_, new_n_n50_,
    new_n__1214_m__, new_n_n73_, new_n__42_m__, new_n_n58_, new_n_n53_,
    new_n_n49_, new_n_n74_, new_n_n63_, new_n_n59_, new_n_n52_,
    new_n__44_m__inv_, new_n_n0_, new_n_n75_, new_n_n43_, new_n_n32_,
    new_n_n21_, new_n_n10_, new_n_n76_, new_n_n42_, new_n_n33_, new_n_n20_,
    new_n_n11_, new_n_n41_, new_n_n30_, new_n_n23_, new_n_n12_, new_n_n40_,
    new_n_n31_, new_n_n22_, new_n_n13_, new_n_n57_, new_n__90_m__,
    new_n__226_m__, new_n_n36_, new_n_n25_, new_n_n14_, new_n_n56_,
    new_n__89_m__, new_n__873_m__, new_n_n37_, new_n_n24_, new_n_n15_,
    new_n_n67_, new_n_n61_, new_n_n45_, new_n_n34_, new_n_n27_, new_n_n16_,
    new_n_n66_, new_n_n62_, new_n_n44_, new_n_n35_, new_n_n26_, new_n_n17_,
    new_n_n68_, new_nc2g5_, new_ntimot_, new_n_n55_, new_n__2087_m__,
    new_n_n29_, new_n_n18_, new_n_n69_, new_n__260_m__, new_n_n60_,
    new_n_n54_, new_n__254_m__inv_, new_n_n28_, new_n_n19_, new_n_n70_,
    new_n__199_m__inv_, new_n__58_m__inv_, new_n__894_m__, new_n__80_m__,
    new_n_n47_, new_n_n38_, new_n_n71_, new_n_n65_, new_n__886_m__,
    new_nc1g3_, new_n__99_m__, new_n_n46_, new_n_n39_;
  assign pbull2_p = new_nbull2_p_;
  assign new_ndel1_ = pdel1;
  assign pend_p = new_nend_p_;
  assign pbull3_p = new_nbull3_p_;
  assign porwd_f = new_norwd_f_;
  assign pbull4_p = new_nbull4_p_;
  assign ppluto3_p = new_npluto3_p_;
  assign pwatch_p = new_nwatch_p_;
  assign pbull5_p = new_nbull5_p_;
  assign new_nratr_ = pratr;
  assign new_nbull1_ = pbull1;
  assign pbull6_p = new_nbull6_p_;
  assign ppluto5_p = new_npluto5_p_;
  assign ppy_p = new_npy_p_;
  assign new_nbull0_ = pbull0;
  assign new_nwatch_ = pwatch;
  assign new_novacc_ = povacc;
  assign new_nverr_n_ = pverr_n;
  assign ppluto4_p = new_npluto4_p_;
  assign plsd_p = new_nlsd_p_;
  assign pvlenesr_p = new_nvlenesr_p_;
  assign new_norwd_n_ = porwd_n;
  assign pfbi_p = new_nfbi_p_;
  assign new_nvlenesr_ = pvlenesr;
  assign pstar1_p = new_nstar1_p_;
  assign pvsumesr_p = new_nvsumesr_p_;
  assign paccrpy_p = new_naccrpy_p_;
  assign pkbg_f = new_nkbg_f_;
  assign pmarssr_p = new_nmarssr_p_;
  assign new_nmmerr_ = pmmerr;
  assign pstar0_p = new_nstar0_p_;
  assign new_naccrpy_ = paccrpy;
  assign pstar3_p = new_nstar3_p_;
  assign pdel1_p = new_ndel1_p_;
  assign pstar2_p = new_nstar2_p_;
  assign new_nvacc_ = pvacc;
  assign new_ncat4_ = pcat4;
  assign new_nvst1_ = pvst1;
  assign new_ncapsd_ = pcapsd;
  assign new_ncat3_ = pcat3;
  assign new_ncat2_ = pcat2;
  assign pvst0_p = new_nvst0_p_;
  assign new_ncat1_ = pcat1;
  assign new_nlsd_ = plsd;
  assign new_nvst0_ = pvst0;
  assign new_ncat0_ = pcat0;
  assign pcomppar_p = new_ncomppar_p_;
  assign new_nibt2_ = pibt2;
  assign new_nkbg_n_ = pkbg_n;
  assign powl_f = new_nowl_f_;
  assign new_nmarssr_ = pmarssr;
  assign psdo = new_nvst0_;
  assign new_nend_ = pend;
  assign pvst1_p = new_nvst1_p_;
  assign new_nvsumesr_ = pvsumesr;
  assign new_nbull5_ = pbull5;
  assign ppluto1_p = new_npluto1_p_;
  assign new_npluto4_ = ppluto4;
  assign new_nstar2_ = pstar2;
  assign new_nbull4_ = pbull4;
  assign new_npluto5_ = ppluto5;
  assign new_npy_ = ppy;
  assign new_nstar3_ = pstar3;
  assign new_nbull3_ = pbull3;
  assign new_ncomppar_ = pcomppar;
  assign new_nibt1_ = pibt1;
  assign pratr_p = new_nratr_p_;
  assign new_nstar0_ = pstar0;
  assign new_nbull2_ = pbull2;
  assign new_nibt0_ = pibt0;
  assign ppluto0_p = new_npluto0_p_;
  assign new_nstar1_ = pstar1;
  assign new_npluto0_ = ppluto0;
  assign new_nfbi_ = pfbi;
  assign povacc_p = new_novacc_p_;
  assign new_nowl_n_ = powl_n;
  assign new_npluto1_ = ppluto1;
  assign ppluto2_p = new_npluto2_p_;
  assign pbull0_p = new_nbull0_p_;
  assign new_niclr_ = piclr;
  assign new_npluto2_ = ppluto2;
  assign pverr_f = new_nverr_f_;
  assign pbull1_p = new_nbull1_p_;
  assign new_nbull6_ = pbull6;
  assign new_ncat5_ = pcat5;
  assign new_npluto3_ = ppluto3;
  assign new_naccrpy_p_ = new_n_n121_ | new_n_n146_;
  assign new_n_n119_ = new_n_n40_ & new_n_n9_ & new_n_n35_;
  assign new_n_n111_ = new_n_n2_ & new_nkbg_n_;
  assign new_nvst1_p_ = new_n_n102_ | new_n_n103_;
  assign new_nstar2_p_ = new_n_n92_ | new_n_n94_ | new_n_n93_ | new_n_n95_;
  assign new_n_n87_ = new_n_n20_ & new_n_n42_;
  assign new_nbull4_p_ = new_n_n79_ | new_n_n78_ | new_n_n77_;
  assign new_n_n147_ = new_nfbi_ & new_n_n6_ & new_n_n35_ & new_n_n14_;
  assign new_n_n118_ = new_n_n37_ & new_n_n9_ & new_n_n35_;
  assign new_nkbg_f_ = new_n_n111_ | new_n_n110_ | new_n_n109_;
  assign new_n_n103_ = new_n__89_m__ & new_nvst1_;
  assign new_n_n96_ = new_nstar0_ & new_n_n37_ & new_n_n13_;
  assign new_n_n86_ = new_nbull0_ & new_nowl_n_ & new_n_n41_;
  assign new_n_n80_ = new_nowl_n_ & new_n_n16_ & new_n_n45_;
  assign new_n_n148_ = new_nc2g5_ & new_nlsd_ & new_nowl_n_;
  assign new_npluto3_p_ = new_n_n130_ | new_n_n131_;
  assign new_n_n125_ = new_n_n41_ & new_n_n19_ & new_nkbg_n_ & new_n_n34_;
  assign new_n_n102_ = new_n__90_m__ & new_npy_;
  assign new_n_n94_ = new_n_n6_ & new_n__99_m__;
  assign new_n_n88_ = new_nstar2_ & new_n_n9_ & new_n__80_m__ & new_n_n14_;
  assign new_n_n81_ = new_nowl_n_ & new_nbull3_ & new_n__226_m__;
  assign new_n_n149_ = new_n_n14_ & new_nlsd_ & new_nowl_n_;
  assign new_n_n131_ = new_nowl_n_ & new_npluto3_;
  assign new_nowl_f_ = new_n_n124_ | new_n_n125_;
  assign new_nstar0_p_ = new_n_n100_ | new_n_n101_;
  assign new_n_n95_ = new_n_n7_ & new_nstar2_;
  assign new_nbull0_p_ = new_n_n86_ | new_n_n87_;
  assign new_nbull3_p_ = new_n_n80_ | new_n_n81_;
  assign new_n_n144_ = new_nverr_n_ & new_n_n2_ & new_n_n0_;
  assign new_npluto0_p_ = new_n_n136_ | new_n_n137_;
  assign new_n_n101_ = new_n_n9_ & new_n_n5_;
  assign new_n_n92_ = new_n_n8_ & new_n__80_m__ & new_n_n13_;
  assign new_n_n84_ = new_n_n43_ & new_nbull0_ & new_n_n20_;
  assign new_nbull5_p_ = new_n_n73_ | new_n_n75_ | new_n_n74_ | new_n_n76_;
  assign new_n_n9_ = ~new_n__254_m__inv_;
  assign new_n_n145_ = new_nverr_n_ & new_n_n41_ & new_n_n2_;
  assign new_n_n143_ = new_nverr_n_ & new_n__42_m__ & new_n_n0_;
  assign new_n_n138_ = new_n_n22_ & new_nvst1_;
  assign new_n_n100_ = new_n_n7_ & new_nstar0_;
  assign new_n_n93_ = new_n__2087_m__ & new_nstar2_;
  assign new_nbull2_p_ = new_n_n82_ | new_n_n83_;
  assign new_n_n77_ = new_nbull4_ & new_nowl_n_ & new_n__226_m__;
  assign new_nverr_f_ = new_n_n143_ | new_n_n145_ | new_n_n144_ | new_n_n109_;
  assign new_nstar1_p_ = new_n_n96_ | new_n_n98_ | new_n_n97_ | new_n_n99_;
  assign new_n_n91_ = new_n_n7_ & new_nstar3_;
  assign new_nbull1_p_ = new_n_n84_ | new_n_n85_;
  assign new_n_n78_ = new_nbull4_ & new_nowl_n_ & new_n_n16_;
  assign new_n_n146_ = new_nowl_n_ & new_naccrpy_;
  assign new_n_n99_ = new_n_n7_ & new_nstar1_;
  assign new_nstar3_p_ = new_n_n88_ | new_n_n90_ | new_n_n89_ | new_n_n91_;
  assign new_n_n85_ = new_n__1214_m__ & new_nbull1_;
  assign new_n_n79_ = new_n__873_m__ & new_n_n10_;
  assign new_nmarssr_p_ = new_n_n59_ | new_n_n141_;
  assign new_n_n135_ = new_nowl_n_ & new_npluto1_;
  assign new_npluto5_p_ = new_n_n126_ | new_n_n127_;
  assign new_n_n121_ = new_n_n13_ & new_n_n2_;
  assign new_n_n112_ = new_n_n1_ & new_nowl_n_ & new_novacc_;
  assign new_nvst0_p_ = new_n_n104_ | new_n_n105_;
  assign new_n_n5_ = ~new_nstar0_;
  assign new_n_n141_ = new_nowl_n_ & new_nmarssr_;
  assign new_npluto1_p_ = new_n_n134_ | new_n_n135_;
  assign new_n_n127_ = new_nowl_n_ & new_npluto5_;
  assign new_nend_p_ = new_n_n121_ | new_n_n22_;
  assign new_novacc_p_ = new_n_n34_ & new_nvacc_;
  assign new_n_n106_ = new_n_n3_ & new_ncomppar_ & new_nowl_n_;
  assign new_n_n6_ = ~new_nc2g5_;
  assign new_nratr_p_ = new_n__886_m__ | new_n_n142_ | new_n_n58_;
  assign new_n_n136_ = new_n_n31_ & new_n__1015_m__ & new_n__894_m__;
  assign new_n_n126_ = new_nibt1_ & new_nibt2_ & new_n__1015_m__ & new_nibt0_;
  assign new_n_n120_ = new_n_n35_ & new_nfbi_;
  assign new_n_n113_ = new_n__99_m__ & new_nstar2_ & new_n__2087_m__ & new_nc2g5_;
  assign new_n_n107_ = new_n_n33_ & new_ncomppar_ & new_nowl_n_;
  assign new_n_n7_ = ~new_n__44_m__inv_;
  assign new_n_n142_ = new_nowl_n_ & new_nratr_;
  assign new_n_n137_ = new_nowl_n_ & new_npluto0_;
  assign new_norwd_f_ = new_n_n12_ | new_n_n41_;
  assign new_nfbi_p_ = new_n_n117_ | new_n_n116_ | new_n_n119_ | new_n_n118_ | new_n_n115_ | new_n_n114_ | new_n_n120_ | new_n_n113_;
  assign new_nwatch_p_ = new_n_n112_ | new_n_n20_;
  assign new_n_n108_ = new_ndel1_ & new_n_n21_ & new_n_n13_;
  assign new_n_n8_ = ~new_nstar2_;
  assign new_n_n150_ = new_n_n33_ & new_nlsd_ & new_nowl_n_;
  assign new_nvsumesr_p_ = new_n_n138_ | new_n_n139_;
  assign new_n_n132_ = new_n_n30_ & new_nibt2_ & new_n__1015_m__ & new_n_n31_;
  assign new_n_n130_ = new_n_n30_ & new_nibt2_ & new_n__1015_m__ & new_nibt0_;
  assign new_npy_p_ = new_n_n122_ | new_n_n123_;
  assign new_n_n115_ = new_n_n37_ & new_nc2g5_ & new_n_n13_;
  assign new_ncomppar_p_ = new_n_n108_ | new_n_n107_ | new_n_n106_;
  assign new_n_n90_ = new_n__2087_m__ & new_nstar3_;
  assign new_n_n82_ = new_nbull1_ & new_nbull0_ & new_n_n20_ & new_n_n44_;
  assign new_n_n1_ = ~new_nvacc_;
  assign new_nlsd_p_ = new_n_n147_ | new_n_n149_ | new_n_n148_ | new_n_n150_;
  assign new_n_n139_ = new_nowl_n_ & new_nvsumesr_;
  assign new_n_n133_ = new_nowl_n_ & new_npluto2_;
  assign new_npluto4_p_ = new_n_n128_ | new_n_n129_;
  assign new_n_n124_ = new_n_n0_ & new_n_n19_ & new_nkbg_n_ & new_n_n34_;
  assign new_n_n114_ = new_nfbi_ & new_nstar2_ & new_n__2087_m__ & new_nc2g5_;
  assign new_ndel1_p_ = new_n_n34_ & new_ncapsd_;
  assign new_n_n89_ = new_nowl_n_ & new_n_n8_ & new_nstar3_;
  assign new_n_n83_ = new_n__1214_m__ & new_nbull2_;
  assign new_n_n2_ = ~new_n__199_m__inv_;
  assign new_nvlenesr_p_ = new_n_n56_ | new_n_n140_;
  assign new_npluto2_p_ = new_n_n132_ | new_n_n133_;
  assign new_n_n129_ = new_nowl_n_ & new_npluto4_;
  assign new_n_n122_ = new_n__90_m__ & new_ndel1_;
  assign new_n_n117_ = new_n_n40_ & new_nc2g5_ & new_n_n13_;
  assign new_n_n109_ = new_n__219_m__ & new_n_n38_;
  assign new_n_n105_ = new_n__89_m__ & new_nvst0_;
  assign new_n_n97_ = new_n_n5_ & new_nstar1_ & new_n__2087_m__;
  assign new_n_n3_ = ~new_ndel1_;
  assign new_n_n140_ = new_nowl_n_ & new_nvlenesr_;
  assign new_n_n134_ = new_nibt0_ & new_n__1015_m__ & new_n__894_m__;
  assign new_n_n128_ = new_nibt1_ & new_nibt2_ & new_n__1015_m__ & new_n_n31_;
  assign new_n_n123_ = new_n__89_m__ & new_npy_;
  assign new_n_n116_ = new_nfbi_ & new_nc2g5_ & new_n_n13_;
  assign new_n_n110_ = new_n__42_m__ & new_nkbg_n_;
  assign new_n_n104_ = new_n__90_m__ & new_nvst1_;
  assign new_n_n98_ = new_nstar0_ & new_n_n4_ & new_n__99_m__;
  assign new_n_n4_ = ~new_nstar1_;
  assign new_n_n72_ = new_n__1214_m__ & new_nbull6_;
  assign new_n_n64_ = new_nc2g5_ & new_n_n13_;
  assign new_n__1015_m__ = new_n_n59_ | new_n_n57_ | new_n_n56_ | new_n_n58_ | new_n__886_m__;
  assign new_n_n51_ = new_n_n29_ & new_n_n30_ & new_nibt2_ & new_nibt0_;
  assign new_n_n48_ = new_n_n42_ & new_nowl_n_;
  assign new_nbull6_p_ = new_n_n69_ | new_n_n68_ | new_n_n71_ | new_n_n70_ | new_n_n66_ | new_n_n72_ | new_n_n67_;
  assign new_n__219_m__ = new_n_n33_ | new_n_n38_;
  assign new_nc29g7_ = new_n_n41_ | new_n_n38_;
  assign new_n_n50_ = new_n_n32_ & new_n_n30_ & new_nibt2_ & new_n_n31_;
  assign new_n__1214_m__ = new_n_n48_ | new_n_n47_ | new_n_n46_;
  assign new_n_n73_ = new_nbull5_ & new_nowl_n_ & new_n__226_m__;
  assign new_n__42_m__ = new_n_n60_ | new_n_n62_ | new_n_n61_ | new_n_n63_;
  assign new_n_n58_ = new_n_n22_ & new_n_n21_;
  assign new_n_n53_ = new_n_n27_ & new_nibt1_ & new_nibt2_ & new_nibt0_;
  assign new_n_n49_ = new_n_n39_ & new_n_n40_;
  assign new_n_n74_ = new_nbull5_ & new_nowl_n_ & new_n_n16_;
  assign new_n_n63_ = new_n_n39_ & new_n_n14_;
  assign new_n_n59_ = new_ntimot_ & new_n_n20_;
  assign new_n_n52_ = new_n_n28_ & new_nibt1_ & new_nibt2_ & new_n_n31_;
  assign new_n__44_m__inv_ = new_n_n38_ | new_nfbi_ | new_n_n49_;
  assign new_n_n0_ = ~new_ntimot_;
  assign new_n_n75_ = new_n_n15_ & new_nbull4_ & new_n__873_m__;
  assign new_n_n43_ = ~new_nbull1_;
  assign new_n_n32_ = ~new_ncat2_;
  assign new_n_n21_ = ~new_ncomppar_;
  assign new_n_n10_ = ~new_nbull4_;
  assign new_n_n76_ = new_nbull4_p_ & new_nbull5_;
  assign new_n_n42_ = ~new_nbull0_;
  assign new_n_n33_ = ~new_nfbi_;
  assign new_n_n20_ = ~new_nc29g7_;
  assign new_n_n11_ = ~new_nbull6_;
  assign new_n_n41_ = ~new_nwatch_;
  assign new_n_n30_ = ~new_nibt1_;
  assign new_n_n23_ = ~new_nkbg_n_;
  assign new_n_n12_ = ~new_nc1g3_;
  assign new_n_n40_ = ~new_norwd_n_;
  assign new_n_n31_ = ~new_nibt0_;
  assign new_n_n22_ = ~new_n__58_m__inv_;
  assign new_n_n13_ = ~new_n__219_m__;
  assign new_n_n57_ = new_nvst1_ & new_n_n22_;
  assign new_n__90_m__ = new_nfbi_ & new_n_n34_;
  assign new_n__226_m__ = new_n_n44_ | new_n_n42_ | new_n_n43_ | new_n_n41_;
  assign new_n_n36_ = ~new_n__99_m__;
  assign new_n_n25_ = ~new_ncat1_;
  assign new_n_n14_ = ~new_nstar3_;
  assign new_n_n56_ = new_n_n23_ & new_nowl_n_;
  assign new_n__89_m__ = new_n_n33_ & new_n_n34_;
  assign new_n__873_m__ = new_nowl_n_ & new_nbull3_ & new_n_n45_;
  assign new_n_n37_ = ~new_n__80_m__;
  assign new_n_n24_ = ~new_nibt2_;
  assign new_n_n15_ = ~new_nbull5_;
  assign new_n_n67_ = new_nbull4_ & new_n_n11_ & new_n__873_m__ & new_nbull5_;
  assign new_n_n61_ = new_n_n14_ & new_nwatch_ & new_n_n25_ & new_n_n26_ & new_n__894_m__;
  assign new_n_n45_ = ~new_n__226_m__;
  assign new_n_n34_ = ~new_niclr_;
  assign new_n_n27_ = ~new_ncat5_;
  assign new_n_n16_ = ~new_nbull3_;
  assign new_n_n66_ = new_nbull3_ & new_nbull5_ & new_nbull4_ & new_n__1214_m__ & new_n_n45_;
  assign new_n_n62_ = new_nc2g5_ & new_n_n39_;
  assign new_n_n44_ = ~new_nbull2_;
  assign new_n_n35_ = ~new_n__260_m__;
  assign new_n_n26_ = ~new_ncat0_;
  assign new_n_n17_ = ~new_nvst0_;
  assign new_n_n68_ = new_n_n15_ & new_nbull6_ & new_nowl_n_;
  assign new_nc2g5_ = new_n_n37_ | new_nstar2_;
  assign new_ntimot_ = new_n_n44_ & new_nbull1_ & new_n_n42_ & new_nbull4_ & new_n_n16_ & new_n_n15_ & new_nbull6_;
  assign new_n_n55_ = new_n_n25_ & new_nibt0_ & new_n__894_m__;
  assign new_n__2087_m__ = new_n_n37_ & new_nowl_n_;
  assign new_n_n29_ = ~new_ncat3_;
  assign new_n_n18_ = ~new_nmmerr_;
  assign new_n_n69_ = new_n_n10_ & new_nbull6_ & new_nowl_n_;
  assign new_n__260_m__ = new_nc29g7_ | new_n_n12_;
  assign new_n_n60_ = new_nc2g5_ & new_nwatch_ & new_n_n25_ & new_n_n26_ & new_n__894_m__;
  assign new_n_n54_ = new_n_n31_ & new_n__894_m__ & new_n_n26_;
  assign new_n__254_m__inv_ = new_n__219_m__ & new_n_n36_;
  assign new_n_n28_ = ~new_ncat4_;
  assign new_n_n19_ = ~new_nend_;
  assign new_n_n70_ = new_n_n16_ & new_nbull6_ & new_nowl_n_;
  assign new_n__199_m__inv_ = new_n_n64_ | new_n_n65_;
  assign new_n__58_m__inv_ = new_n_n19_ | new_n_n38_;
  assign new_n__894_m__ = new_n_n24_ & new_nibt1_;
  assign new_n__80_m__ = new_nstar1_ & new_nstar0_;
  assign new_n_n47_ = new_n_n43_ & new_nowl_n_;
  assign new_n_n38_ = ~new_nowl_n_;
  assign new_n_n71_ = new_n_n44_ & new_nbull6_ & new_nowl_n_;
  assign new_n_n65_ = new_n_n13_ & new_n_n39_;
  assign new_n__886_m__ = new_n_n18_ & new_n_n17_ & new_n_n22_;
  assign new_nc1g3_ = new_n_n54_ | new_n_n52_ | new_n_n51_ | new_n_n50_ | new_n_n53_ | new_n_n55_;
  assign new_n__99_m__ = new_n_n35_ & new_n_n40_;
  assign new_n_n46_ = new_n_n41_ & new_nowl_n_;
  assign new_n_n39_ = ~new_norwd_f_;
endmodule


