// Benchmark "top" written by ABC on Fri Mar 31 12:12:53 2023

module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0,
    px, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0, pb, pr0,
    pc, ps0, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po,
    pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pg2, pd2, pg1, pe2, pf1,
    pi1, pj2, ph1, pk2, ph2, pk1, pi2, pj1, pm1, pl1, pl2, po1, pn1, pq1,
    pp1, ps1, pr1, pt0, pu1, pt1, pu0, pv0, pw1, pv1, pw0, px0, py1, px1,
    py0, pz0, pz1  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0,
    pw, ph0, px, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0,
    pb, pr0, pc, ps0, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po;
  output pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pg2, pd2, pg1, pe2, pf1,
    pi1, pj2, ph1, pk2, ph2, pk1, pi2, pj1, pm1, pl1, pl2, po1, pn1, pq1,
    pp1, ps1, pr1, pt0, pu1, pt1, pu0, pv0, pw1, pv1, pw0, px0, py1, px1,
    py0, pz0, pz1;
  wire new_np_, new_na0_, new_nq_, new_nb0_, new_nr_, new_nc0_, new_ns_,
    new_nd0_, new_nt_, new_ne0_, new_nu_, new_nf0_, new_nv_, new_ng0_,
    new_nw_, new_nh0_, new_nx_, new_ni0_, new_ny_, new_nj0_, new_nz_,
    new_nk0_, new_nl0_, new_nm0_, new_nn0_, new_no0_, new_np0_, new_na_,
    new_nq0_, new_nb_, new_nr0_, new_nc_, new_ns0_, new_nd_, new_ne_,
    new_nf_, new_ng_, new_nh_, new_ni_, new_nj_, new_nk_, new_nl_, new_nm_,
    new_nn_, new_no_, new_nd5_, new_nc2_, new_n_n62_, new_n_n51_, new_ni2_,
    new_ng6_, new_nr6_, new_nj8_, new_nu8_, new_nf9_, new_nq9_, new_nb10_,
    new_nm10_, new_nh1_, new_nd2_, new_n_n63_, new_n_n50_, new_nh2_,
    new_nh6_, new_nq6_, new_nk8_, new_nt8_, new_ng9_, new_np9_, new_nc10_,
    new_nl10_, new_ni1_, new_nt1_, new_n_n64_, new_n_n49_, new_nx5_,
    new_ne6_, new_np6_, new_np7_, new_na8_, new_nh9_, new_ns9_, new_nz9_,
    new_nk10_, new_nj1_, new_ns1_, new_nb2_, new_n_n48_, new_nk2_,
    new_nf6_, new_no6_, new_nq7_, new_nz7_, new_ni9_, new_nr9_, new_na10_,
    new_nj10_, new_nz0_, new_n_n47_, new_nz5_, new_nk6_, new_nv6_,
    new_ng7_, new_nj9_, new_nu9_, new_nf10_, new_nq10_, new_n_n9_,
    new_ny0_, new_n_n46_, new_ny5_, new_nu6_, new_nw6_, new_nf7_, new_nk9_,
    new_nt9_, new_ng10_, new_np10_, new_nx0_, new_n_n45_, new_ni6_,
    new_nt6_, new_nl9_, new_nw9_, new_nd10_, new_no10_, new_na6_, new_nj6_,
    new_ns6_, new_nm9_, new_nv9_, new_ne10_, new_nn10_, new_nd1_, new_no1_,
    new_nz1_, new_n_n65_, new_nz6_, new_nk7_, new_nv7_, new_ng8_, new_nr8_,
    new_nc9_, new_n_n5_, new_nj2_, new_nc1_, new_np1_, new_ny1_,
    new_n_n55_, new_na7_, new_nj7_, new_nw7_, new_nf8_, new_ns8_, new_nb9_,
    new_n_n6_, new_nb1_, new_nq1_, new_n_n67_, new_n_n56_, new_nx6_,
    new_ni7_, new_nx7_, new_ni8_, new_np8_, new_na9_, new_n_n7_, new_na1_,
    new_na2_, new_n_n66_, new_n_n57_, new_ny6_, new_nh7_, new_ny7_,
    new_nh8_, new_nq8_, new_nz8_, new_n_n8_, new_nw0_, new_nk1_, new_nv1_,
    new_nf2_, new_n_n58_, new_n_n44_, new_nc6_, new_nn6_, new_nd7_,
    new_no7_, new_nr7_, new_nc8_, new_nn8_, new_ny8_, new_nx9_, new_ni10_,
    new_n_n1_, new_ng1_, new_nl1_, new_nu1_, new_n_n68_, new_n_n59_,
    new_n_n54_, new_nd6_, new_nm6_, new_ne7_, new_nn7_, new_ns7_, new_nb8_,
    new_no8_, new_nx8_, new_ny9_, new_nh10_, new_n_n2_, new_nt0_, new_nf1_,
    new_nm1_, new_nx1_, new_ne2_, new_n_n60_, new_n_n53_, new_ng2_,
    new_nl6_, new_nb7_, new_nm7_, new_nt7_, new_ne8_, new_nl8_, new_nw8_,
    new_nd9_, new_no9_, new_n_n3_, new_nu0_, new_ne1_, new_nn1_, new_nw1_,
    new_n_n69_, new_n_n61_, new_n_n52_, new_n_n43_, new_nb6_, new_nc7_,
    new_nl7_, new_nu7_, new_nd8_, new_nm8_, new_nv8_, new_ne9_, new_nn9_,
    new_n_n4_, new_nw10_, new_nh11_, new_ns11_, new_nd12_, new_no12_,
    new_nv10_, new_ni11_, new_nr11_, new_ne12_, new_nn12_, new_nu10_,
    new_nj11_, new_nu11_, new_nb12_, new_nm12_, new_nt10_, new_nk11_,
    new_nt11_, new_nc12_, new_nl12_, new_n_n0_, new_ns10_, new_nv12_,
    new_n_n32_, new_n_n21_, new_n_n10_, new_nr10_, new_n_n42_, new_n_n33_,
    new_n_n20_, new_n_n11_, new_n_n41_, new_n_n30_, new_n_n23_, new_n_n12_,
    new_n_n40_, new_n_n31_, new_n_n22_, new_n_n13_, new_nv11_, new_ng12_,
    new_nr12_, new_n_n36_, new_n_n25_, new_n_n14_, new_nw11_, new_nf12_,
    new_ns12_, new_n_n37_, new_n_n24_, new_n_n15_, new_nb11_, new_nm11_,
    new_nt12_, new_n_n34_, new_n_n27_, new_n_n16_, new_nc11_, new_nl11_,
    new_nu12_, new_n_n35_, new_n_n26_, new_n_n17_, new_na11_, new_nd11_,
    new_no11_, new_nz11_, new_nk12_, new_n_n29_, new_n_n18_, new_nz10_,
    new_ne11_, new_nn11_, new_na12_, new_nj12_, new_n_n28_, new_n_n19_,
    new_ny10_, new_nf11_, new_nq11_, new_nx11_, new_ni12_, new_np12_,
    new_n_n38_, new_nx10_, new_ng11_, new_np11_, new_ny11_, new_nh12_,
    new_nq12_, new_n_n39_;
  assign pa1 = new_na1_;
  assign pb2 = new_nb2_;
  assign new_np_ = pp;
  assign new_na0_ = pa0;
  assign pc2 = new_nc2_;
  assign new_nq_ = pq;
  assign new_nb0_ = pb0;
  assign pc1 = new_nc1_;
  assign new_nr_ = pr;
  assign pa2 = new_na2_;
  assign pb1 = new_nb1_;
  assign new_nc0_ = pc0;
  assign new_ns_ = ps;
  assign new_nd0_ = pd0;
  assign pe1 = new_ne1_;
  assign pf2 = new_nf2_;
  assign new_nt_ = pt;
  assign pd1 = new_nd1_;
  assign new_ne0_ = pe0;
  assign pg2 = new_ng2_;
  assign new_nu_ = pu;
  assign pd2 = new_nd2_;
  assign new_nf0_ = pf0;
  assign pg1 = new_ng1_;
  assign new_nv_ = pv;
  assign pe2 = new_ne2_;
  assign pf1 = new_nf1_;
  assign new_ng0_ = pg0;
  assign new_nw_ = pw;
  assign new_nh0_ = ph0;
  assign pi1 = new_ni1_;
  assign pj2 = new_nj2_;
  assign new_nx_ = px;
  assign ph1 = new_nh1_;
  assign new_ni0_ = pi0;
  assign pk2 = new_nk2_;
  assign new_ny_ = py;
  assign ph2 = new_nh2_;
  assign new_nj0_ = pj0;
  assign pk1 = new_nk1_;
  assign new_nz_ = pz;
  assign pi2 = new_ni2_;
  assign pj1 = new_nj1_;
  assign new_nk0_ = pk0;
  assign new_nl0_ = pl0;
  assign pm1 = new_nm1_;
  assign pl1 = new_nl1_;
  assign new_nm0_ = pm0;
  assign pl2 = new_nd5_;
  assign new_nn0_ = pn0;
  assign po1 = new_no1_;
  assign pn1 = new_nn1_;
  assign new_no0_ = po0;
  assign new_np0_ = pp0;
  assign pq1 = new_nq1_;
  assign new_na_ = pa;
  assign pp1 = new_np1_;
  assign new_nq0_ = pq0;
  assign new_nb_ = pb;
  assign new_nr0_ = pr0;
  assign ps1 = new_ns1_;
  assign new_nc_ = pc;
  assign pr1 = new_nd5_;
  assign new_ns0_ = ps0;
  assign new_nd_ = pd;
  assign pt0 = new_nt0_;
  assign pu1 = new_nu1_;
  assign new_ne_ = pe;
  assign pt1 = new_nt1_;
  assign pu0 = new_nu0_;
  assign new_nf_ = pf;
  assign pv0 = new_nj2_;
  assign pw1 = new_nw1_;
  assign new_ng_ = pg;
  assign pv1 = new_nv1_;
  assign pw0 = new_nw0_;
  assign new_nh_ = ph;
  assign px0 = new_nx0_;
  assign py1 = new_ny1_;
  assign new_ni_ = pi;
  assign px1 = new_nx1_;
  assign py0 = new_ny0_;
  assign new_nj_ = pj;
  assign pz0 = new_nz0_;
  assign new_nk_ = pk;
  assign pz1 = new_nz1_;
  assign new_nl_ = pl;
  assign new_nm_ = pm;
  assign new_nn_ = pn;
  assign new_no_ = po;
  assign new_nd5_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nw_;
  assign new_nc2_ = new_nd9_ | new_ne9_ | new_nh9_ | new_ni9_ | new_nb6_ | new_no9_ | new_nh8_ | new_nf8_ | new_nc6_ | new_nk8_ | new_ne6_ | new_nj8_ | new_np6_ | new_nx10_ | new_nm6_ | new_nh6_ | new_np9_ | new_no8_ | new_nk6_ | new_nz10_ | new_nn7_ | new_nl8_ | new_nv10_ | new_nw11_ | new_nn6_ | new_nt11_ | new_ne12_ | new_ns6_ | new_nj12_ | new_nf10_ | new_nq8_ | new_nz11_ | new_nd11_ | new_nv12_ | new_na6_ | new_nq6_ | new_nf11_ | new_ny9_ | new_no12_ | new_nx11_ | new_nz5_ | new_nq12_ | new_ni2_ | new_nd12_ | new_na11_ | new_nu7_ | new_ns11_ | new_nc11_ | new_no6_ | new_nr11_ | new_nc12_ | new_nd8_ | new_nx9_ | new_nw10_ | new_no11_ | new_nn11_ | new_np11_ | new_nl10_ | new_nw6_ | new_nh12_ | new_nk10_ | new_nm12_ | new_ng11_ | new_ng10_ | new_nv6_ | new_nt10_ | new_nu6_ | new_nk12_ | new_na9_ | new_nw8_ | new_nx8_ | new_nb9_ | new_nc9_;
  assign new_n_n62_ = new_n_n29_ & new_n_n38_ & new_nz_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nd0_;
  assign new_n_n51_ = new_n_n38_ & new_nd0_ & new_na0_ & new_n_n29_ & new_n_n36_ & new_ns_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_n_n39_;
  assign new_ni2_ = new_nv_ & new_nu_ & new_n_n39_ & new_nw_ & new_n_n37_ & new_ne0_ & new_na_ & new_n_n27_ & new_n_n42_ & new_n_n41_ & new_nt_;
  assign new_ng6_ = new_ne0_ & new_nd0_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nz_;
  assign new_nr6_ = new_nc0_ & new_na0_ & new_n_n38_ & new_n_n37_ & new_nr_ & new_n_n35_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_nj8_ = new_n_n30_ & new_n_n40_ & new_nd0_ & new_nc0_ & new_n_n38_ & new_n_n29_ & new_ns_ & new_n_n18_ & new_nt_ & new_nu_;
  assign new_nu8_ = new_n_n38_ & new_n_n37_ & new_nn_ & new_nv_ & new_n_n20_ & new_n_n30_ & new_n_n39_;
  assign new_nf9_ = new_ne0_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_na0_;
  assign new_nq9_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_n_n28_ & new_nt_ & new_n_n41_ & new_nv_ & new_nz_;
  assign new_nb10_ = new_ne0_ & new_ns_ & new_nu_ & new_nt_ & new_nv_ & new_nd0_;
  assign new_nm10_ = new_nd0_ & new_n_n39_ & new_ne0_ & new_ns_ & new_nu_ & new_n_n35_ & new_nv_ & new_nw_;
  assign new_nh1_ = new_nh11_ | new_nn12_ | new_ne11_ | new_ni12_ | new_nt9_ | new_ni8_ | new_nr11_ | new_no12_ | new_no1_ | new_nh8_ | new_nn1_ | new_nx7_ | new_nr6_ | new_nv7_ | new_nc8_ | new_nz7_ | new_no11_ | new_nd6_ | new_ny5_ | new_nt7_ | new_ng6_ | new_nj6_ | new_nf9_ | new_nr7_ | new_nz9_ | new_na11_ | new_np9_ | new_nt6_;
  assign new_nd2_ = new_ni9_ | new_nm9_ | new_ne9_ | new_nl6_ | new_nw9_ | new_nn9_ | new_np8_ | new_nx10_ | new_no6_ | new_nv12_ | new_nj11_ | new_nb6_ | new_nd6_ | new_nd11_ | new_ng10_ | new_ns11_ | new_nc7_ | new_nq8_ | new_ng11_ | new_nm8_ | new_nr12_ | new_nj8_ | new_nq12_ | new_ny10_ | new_na10_ | new_nh8_ | new_nv11_ | new_no10_ | new_ny9_ | new_nu6_ | new_na11_ | new_nk6_ | new_nn10_ | new_ng8_ | new_nd12_ | new_nc8_ | new_nr6_ | new_np6_ | new_ns8_ | new_nr7_ | new_nz1_ | new_nx8_ | new_nt8_ | new_nv8_ | new_nl10_ | new_ne6_ | new_nx9_ | new_nu7_ | new_nt11_ | new_ni10_;
  assign new_n_n63_ = new_n_n29_ & new_ne0_ & new_nz_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_n_n37_;
  assign new_n_n50_ = new_n_n38_ & new_nd0_ & new_n_n30_ & new_n_n29_ & new_n_n18_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_nc0_;
  assign new_nh2_ = new_no8_ | new_nv9_ | new_nt12_ | new_nc10_ | new_nd10_ | new_np10_ | new_nx5_;
  assign new_nh6_ = new_n_n37_ & new_nz_ & new_ne0_ & new_nk_ & new_nt_ & new_ns_ & new_n_n34_ & new_n_n40_;
  assign new_nq6_ = new_na0_ & new_n_n40_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_na_ & new_ns_ & new_n_n26_ & new_n_n35_ & new_nu_;
  assign new_nk8_ = new_nc0_ & new_n_n30_ & new_n_n38_ & new_nd0_ & new_ne_ & new_nt_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_nt8_ = new_n_n39_ & new_n_n30_ & new_n_n38_ & new_n_n37_ & new_n_n20_ & new_n_n35_ & new_ns_ & new_n_n34_ & new_n_n40_;
  assign new_ng9_ = new_n_n37_ & new_ny_ & new_ne0_ & new_n_n29_ & new_n_n35_ & new_n_n41_ & new_nu_ & new_nv_;
  assign new_np9_ = new_n_n39_ & new_nx_ & new_ne0_ & new_n_n37_ & new_nb_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nc10_ = new_nd0_ & new_n_n39_ & new_n_n38_ & new_nd_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_n_n40_;
  assign new_nl10_ = new_nd0_ & new_n_n39_ & new_n_n38_ & new_ns_ & new_nu_ & new_n_n35_ & new_nv_ & new_nw_;
  assign new_ni1_ = new_np9_ | new_ny9_ | new_no9_ | new_nf10_ | new_no6_ | new_ni7_ | new_ng7_ | new_nl7_ | new_nj7_ | new_nu11_ | new_ni10_ | new_ng10_ | new_nm7_ | new_nn7_ | new_nx11_ | new_ni12_ | new_no7_ | new_nj6_ | new_ng6_ | new_nn12_ | new_nd11_ | new_ns7_ | new_nu12_ | new_nd7_ | new_ne8_ | new_nc6_ | new_nq11_ | new_na11_ | new_nf6_ | new_nt12_ | new_nf8_ | new_ny11_ | new_nx10_ | new_ny5_ | new_nu9_ | new_nz11_ | new_nl10_ | new_nm8_ | new_ng12_ | new_nm12_ | new_nc10_ | new_nl12_ | new_nd10_ | new_no8_ | new_nr11_ | new_nw6_ | new_nx9_ | new_nk8_ | new_no1_ | new_nf12_ | new_ng11_ | new_ni8_ | new_ne9_ | new_ni9_ | new_nu8_ | new_nx8_ | new_nr8_ | new_ng8_ | new_nn1_ | new_nk12_;
  assign new_nt1_ = new_ne12_ | new_nc12_ | new_nj12_ | new_np11_;
  assign new_n_n64_ = new_n_n29_ & new_ne0_ & new_na0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_n_n37_;
  assign new_n_n49_ = new_nd0_ & new_n_n39_ & new_n_n29_ & new_n_n38_ & new_n_n42_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_nx5_ = new_nz_ & new_nv_ & new_n_n37_ & new_n_n39_ & new_ne0_ & new_nf_ & new_ns_ & new_nk_ & new_n_n35_ & new_nu_;
  assign new_ne6_ = new_n_n40_ & new_n_n34_ & new_nd0_ & new_nz_ & new_n_n38_ & new_na_ & new_n_n26_ & new_nk_ & new_ns_ & new_nt_;
  assign new_np6_ = new_n_n40_ & new_n_n34_ & new_nd0_ & new_nz_ & new_n_n38_ & new_na_ & new_nl_ & new_nk_ & new_ns_ & new_nt_;
  assign new_np7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_n_n10_ & new_n_n14_ & new_n_n8_ & new_n_n9_ & new_n_n11_ & new_n_n12_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_na8_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_n_n16_ & new_n_n14_ & new_n_n15_ & new_nj_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nh9_ = new_n_n37_ & new_ny_ & new_ne0_ & new_na_ & new_n_n35_ & new_n_n41_ & new_nu_ & new_nv_;
  assign new_ns9_ = new_nd0_ & new_n_n39_ & new_n_n38_ & new_n_n41_ & new_n_n34_ & new_nt_ & new_nv_ & new_nx_;
  assign new_nz9_ = new_nd0_ & new_n_n39_ & new_ne0_ & new_n_n41_ & new_nu_ & new_nt_ & new_nv_ & new_nw_;
  assign new_nk10_ = new_nv_ & new_nu_ & new_n_n39_ & new_nw_ & new_n_n37_ & new_ne0_ & new_na_ & new_n_n27_ & new_n_n42_ & new_ns_ & new_n_n35_;
  assign new_nj1_ = new_nc10_ | new_nx11_ | new_ng11_ | new_nd10_ | new_nq11_ | new_nd5_ | new_nr11_ | new_no11_ | new_na12_ | new_nj6_ | new_nq7_ | new_nk8_ | new_nh6_ | new_ni8_ | new_ni12_ | new_nt7_ | new_nc6_ | new_nw6_ | new_nu7_ | new_nh8_ | new_nn12_ | new_ng6_ | new_nv6_ | new_nv7_ | new_ng8_ | new_nu9_ | new_nk12_ | new_ny7_ | new_nr6_ | new_ns12_ | new_nx7_ | new_nm8_ | new_nn1_ | new_np12_ | new_no8_ | new_nr8_ | new_nw7_ | new_na11_ | new_nd11_ | new_nu8_ | new_ne9_ | new_no12_ | new_nq8_ | new_no1_ | new_nt12_ | new_nz7_ | new_ne12_ | new_nn6_ | new_ny5_ | new_nf12_ | new_ne8_ | new_ny6_ | new_nd8_ | new_nd6_;
  assign new_ns1_ = new_nm11_ | new_nd5_ | new_nk11_ | new_nz11_ | new_np11_ | new_ny6_ | new_nc12_ | new_ni6_ | new_nj12_ | new_nw6_ | new_nv10_ | new_nn6_ | new_np12_ | new_nx6_ | new_nb12_ | new_nm12_ | new_nz6_ | new_nv6_ | new_nb7_ | new_ne12_ | new_nq10_ | new_nn7_ | new_nr10_ | new_ns10_ | new_nz8_ | new_nq9_ | new_nu8_ | new_nc6_ | new_ns12_ | new_nh6_;
  assign new_nb2_ = new_nz9_ | new_nh10_ | new_nm10_ | new_ny10_ | new_ni10_ | new_nu11_ | new_ne11_ | new_ns11_ | new_no11_ | new_nw7_ | new_nm8_ | new_nn8_ | new_nj11_ | new_nv7_ | new_nq6_ | new_nt7_ | new_nj8_ | new_nd7_ | new_nl8_ | new_ns6_ | new_nr7_ | new_ng12_ | new_nx11_ | new_nq7_ | new_nb8_ | new_nv11_ | new_nc8_ | new_nr6_ | new_nz7_ | new_nz5_ | new_nr12_ | new_no7_ | new_na6_ | new_no12_ | new_na8_ | new_nf6_ | new_nu12_ | new_nx7_ | new_nd6_ | new_nk12_ | new_nm9_ | new_nm6_ | new_no6_ | new_ny7_ | new_nn9_ | new_nl6_;
  assign new_n_n48_ = new_n_n38_ & new_nd0_ & new_n_n32_ & new_n_n29_ & new_n_n42_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_n_n40_ & new_n_n39_;
  assign new_nk2_ = new_nz11_ | new_nd5_;
  assign new_nf6_ = new_nd0_ & new_n_n39_ & new_ne0_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_na0_;
  assign new_no6_ = new_n_n38_ & new_n_n41_ & new_nv_ & new_nt_ & new_nc0_ & new_nd0_;
  assign new_nq7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_n_n10_ & new_n_n14_ & new_ns0_ & new_n_n9_ & new_n_n11_ & new_n_n12_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nz7_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_n_n16_ & new_nn0_ & new_n_n15_ & new_nj_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_ni9_ = new_n_n38_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_ny_;
  assign new_nr9_ = new_nd0_ & new_n_n39_ & new_n_n38_ & new_n_n41_ & new_n_n34_ & new_nt_ & new_nv_ & new_nw_;
  assign new_na10_ = new_nw_ & new_nv_ & new_n_n37_ & new_nc0_ & new_n_n38_ & new_n_n22_ & new_n_n41_ & new_nq_ & new_nt_ & new_nu_;
  assign new_nj10_ = new_ne0_ & new_n_n37_ & new_ns_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nc0_;
  assign new_nz0_ = new_nk10_ | new_nz10_ | new_ni2_ | new_nc11_ | new_nw10_ | new_ns6_ | new_nt11_ | new_na6_ | new_nk12_ | new_np6_ | new_nd12_ | new_nb6_ | new_nv12_ | new_nk6_ | new_nf11_ | new_nx11_ | new_nq6_ | new_ne6_ | new_nq12_ | new_nj8_ | new_nu6_ | new_ng8_ | new_nc9_ | new_nd9_ | new_na9_ | new_nb9_ | new_nw8_ | new_nn8_ | new_ns11_ | new_nz5_;
  assign new_n_n47_ = new_ne0_ & new_nd0_ & new_n_n30_ & new_n_n29_ & new_n_n42_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_n_n39_;
  assign new_nz5_ = new_na0_ & new_n_n40_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_na_ & new_ns_ & new_n_n26_ & new_nt_ & new_n_n34_;
  assign new_nk6_ = new_nd0_ & new_nw_ & new_n_n38_ & new_na_ & new_nt_ & new_ns_ & new_n_n34_ & new_n_n40_;
  assign new_nv6_ = new_n_n39_ & new_na0_ & new_ne0_ & new_n_n37_ & new_n_n36_ & new_n_n35_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_ng7_ = new_n_n38_ & new_nd0_ & new_n_n7_ & new_n_n16_ & new_n_n15_ & new_n_n5_ & new_n_n6_ & new_nl0_ & new_n_n4_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_nj9_ = new_ne0_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_ny_;
  assign new_nu9_ = new_nw_ & new_n_n40_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_nc_ & new_n_n41_ & new_n_n32_ & new_nt_ & new_nu_;
  assign new_nf10_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_na_ & new_n_n35_ & new_ns_ & new_n_n34_ & new_nv_;
  assign new_nq10_ = new_ne0_ & new_ns_ & new_n_n34_ & new_n_n35_ & new_n_n40_ & new_nw_;
  assign new_n_n9_ = ~new_nr0_;
  assign new_ny0_ = new_nt10_ | new_nm6_ | new_nf10_ | new_nh9_;
  assign new_n_n46_ = new_ne0_ & new_n_n37_ & new_n_n42_ & new_n_n29_ & new_n_n27_ & new_ns_ & new_nu_ & new_n_n35_ & new_nv_ & new_n_n39_;
  assign new_ny5_ = new_nd0_ & new_nc0_ & new_n_n38_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_na0_;
  assign new_nu6_ = new_na0_ & new_n_n40_ & new_nd0_ & new_n_n39_ & new_n_n38_ & new_na_ & new_ns_ & new_nr_ & new_n_n35_ & new_nu_;
  assign new_nw6_ = new_n_n39_ & new_na0_ & new_ne0_ & new_n_n37_ & new_nr_ & new_n_n35_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_nf7_ = new_n_n38_ & new_nd0_ & new_n_n7_ & new_n_n16_ & new_n_n15_ & new_n_n5_ & new_n_n6_ & new_n_n3_ & new_n_n4_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_nk9_ = new_nw_ & new_nv_ & new_n_n37_ & new_nc0_ & new_n_n38_ & new_nh_ & new_n_n41_ & new_n_n25_ & new_nt_ & new_nu_;
  assign new_nt9_ = new_ne0_ & new_ns_ & new_n_n34_ & new_nt_ & new_nv_ & new_na0_;
  assign new_ng10_ = new_n_n38_ & new_nd0_ & new_ns_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_n_n39_;
  assign new_np10_ = new_n_n39_ & new_n_n24_ & new_ne0_ & new_n_n37_ & new_nf_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_nx0_ = new_nl6_ | new_nn9_ | new_nl11_;
  assign new_n_n45_ = new_ne0_ & new_n_n37_ & new_n_n32_ & new_n_n29_ & new_nc_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nc0_;
  assign new_ni6_ = new_n_n37_ & new_nz_ & new_ne0_ & new_n_n28_ & new_nt_ & new_ns_ & new_n_n34_ & new_n_n40_;
  assign new_nt6_ = new_ne0_ & new_n_n41_ & new_nv_ & new_nt_ & new_nc0_ & new_nd0_;
  assign new_nl9_ = new_ne0_ & new_nz_ & new_nk_ & new_nt_ & new_ns_ & new_n_n34_ & new_nv_;
  assign new_nw9_ = new_nw_ & new_nv_ & new_n_n37_ & new_n_n39_ & new_ne0_ & new_n_n42_ & new_n_n41_ & new_np_ & new_nt_ & new_nu_;
  assign new_nd10_ = new_n_n39_ & new_n_n40_ & new_n_n38_ & new_nd0_ & new_n_n32_ & new_n_n41_ & new_nf_ & new_n_n35_ & new_n_n34_;
  assign new_no10_ = new_nc0_ & new_nv_ & new_n_n23_ & new_ns_ & new_n_n25_ & new_n_n35_ & new_nu_;
  assign new_na6_ = new_na0_ & new_n_n40_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_na_ & new_ns_ & new_nl_ & new_nt_ & new_n_n34_;
  assign new_nj6_ = new_ne0_ & new_nd0_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_ns6_ = new_na0_ & new_n_n40_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_na_ & new_ns_ & new_nl_ & new_n_n35_ & new_nu_;
  assign new_nm9_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_nk_ & new_nt_ & new_n_n41_ & new_nv_ & new_nz_;
  assign new_nv9_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_nf_ & new_nt_ & new_n_n41_ & new_nu_ & new_nv_;
  assign new_ne10_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_n_n29_ & new_n_n35_ & new_ns_ & new_n_n34_ & new_nv_;
  assign new_nn10_ = new_n_n39_ & new_nv_ & new_ne0_ & new_n_n37_ & new_n_n42_ & new_ns_ & new_np_ & new_n_n35_ & new_nu_;
  assign new_nd1_ = new_np9_ | new_no6_ | new_ng10_ | new_nl10_ | new_ny9_ | new_na11_ | new_nx10_ | new_nl12_ | new_nn12_ | new_nv7_ | new_ny5_ | new_nu7_ | new_nf6_ | new_nh11_ | new_ni8_ | new_nr11_ | new_nt7_ | new_ng12_ | new_ng11_ | new_nm8_ | new_ne11_ | new_nq7_ | new_nd8_ | new_ni12_ | new_nd11_ | new_nf8_ | new_nu12_ | new_ny11_ | new_nz7_ | new_ng6_ | new_nd7_ | new_ny7_ | new_nj6_ | new_ne9_ | new_ni9_ | new_no9_ | new_nx7_ | new_nf9_ | new_nx8_ | new_nn1_ | new_nu11_ | new_nw7_ | new_no1_ | new_nx9_;
  assign new_no1_ = new_nd0_ & new_nc0_ & new_n_n38_ & new_ns_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_na0_;
  assign new_nz1_ = new_n_n37_ & new_n_n39_ & new_n_n38_ & new_n_n1_ & new_n_n20_ & new_n_n0_ & new_nv_ & new_n_n30_;
  assign new_n_n65_ = new_n_n38_ & new_nd0_ & new_n_n29_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_nz6_ = new_ne0_ & new_nz_ & new_n_n28_ & new_n_n35_ & new_ns_ & new_n_n34_ & new_n_n40_;
  assign new_nk7_ = new_n_n38_ & new_nd0_ & new_n_n7_ & new_n_n16_ & new_nh0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_nv7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_n_n12_ & new_nn0_ & new_n_n11_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_ng8_ = new_nb0_ & new_n_n40_ & new_n_n38_ & new_n_n37_ & new_na_ & new_ns_ & new_nd_ & new_nt_ & new_nu_;
  assign new_nr8_ = new_no_ & new_n_n39_ & new_n_n30_ & new_n_n37_ & new_n_n38_;
  assign new_nc9_ = new_na0_ & new_nv_ & new_ne0_ & new_n_n37_ & new_na_ & new_n_n41_ & new_n_n26_ & new_n_n35_ & new_nu_;
  assign new_n_n5_ = ~new_nj0_;
  assign new_nj2_ = 1'b0;
  assign new_nc1_ = new_nx11_ | new_nd12_ | new_ng8_;
  assign new_np1_ = new_ni9_ | new_no9_ | new_nf9_ | new_np9_ | new_nj9_ | new_ny6_ | new_ns12_ | new_nj6_ | new_nd8_ | new_nq8_ | new_nx6_ | new_np12_ | new_no8_ | new_nn6_ | new_ne8_ | new_nb7_ | new_nj12_ | new_nm8_ | new_nh6_ | new_ni12_ | new_nf8_ | new_ni6_ | new_nz6_ | new_ng8_ | new_nk8_ | new_ni10_ | new_nr9_ | new_no11_ | new_nv10_ | new_nr6_ | new_nx7_ | new_nf6_ | new_nj10_ | new_nq9_ | new_nu9_ | new_nn12_ | new_ng12_ | new_ny7_ | new_nd6_ | new_np11_ | new_ne11_ | new_no12_ | new_nm12_ | new_no1_ | new_nz7_ | new_ny5_ | new_nc10_ | new_nd11_ | new_nr11_ | new_nk12_ | new_ne12_ | new_nn1_ | new_ny9_ | new_nc8_ | new_nh11_ | new_nr10_ | new_nf12_ | new_nd10_ | new_na12_ | new_nw7_ | new_ni8_ | new_nf10_ | new_nl7_ | new_nb10_ | new_nx10_ | new_nx9_ | new_ny10_ | new_nu7_ | new_nd7_ | new_nz9_ | new_nk7_ | new_nt7_ | new_nc12_ | new_nj7_ | new_ni7_ | new_nr7_ | new_nh7_ | new_ns7_ | new_np7_ | new_nr8_ | new_nz8_ | new_ne9_ | new_no7_ | new_nx8_ | new_nn7_ | new_ny8_ | new_nq7_ | new_ng7_ | new_nm10_ | new_nd5_ | new_ni11_ | new_nc6_ | new_nw6_ | new_na11_ | new_nh10_ | new_nz11_ | new_nk11_ | new_nv7_ | new_nh8_ | new_ng10_ | new_nm7_ | new_nt9_ | new_nb11_ | new_nt12_ | new_ns10_ | new_nt6_ | new_nu11_ | new_ng11_ | new_nu12_ | new_nq11_ | new_nv6_ | new_nx11_ | new_ns9_ | new_ng6_ | new_no6_ | new_nl9_ | new_nl10_;
  assign new_ny1_ = new_nq6_ | new_na6_ | new_nz5_ | new_nj8_ | new_ns6_ | new_ns11_;
  assign new_n_n55_ = new_n_n37_ & new_n_n39_ & new_nx_ & new_ne0_ & new_n_n2_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_na7_ = new_nw_ & new_nv_ & new_n_n37_ & new_nc0_ & new_n_n38_ & new_ni_ & new_n_n41_ & new_nq_ & new_nt_ & new_nu_;
  assign new_nj7_ = new_n_n38_ & new_nd0_ & new_n_n7_ & new_n_n16_ & new_n_n15_ & new_ni0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_nw7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_n_n12_ & new_n_n14_ & new_nq0_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nf8_ = new_ne0_ & new_n_n37_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_nb0_;
  assign new_ns8_ = new_n_n30_ & new_n_n19_ & new_n_n37_ & new_n_n39_ & new_n_n38_ & new_n_n20_ & new_n_n35_ & new_n_n41_ & new_nu_ & new_n_n40_;
  assign new_nb9_ = new_nv_ & new_nu_ & new_n_n37_ & new_nz_ & new_ne0_ & new_na_ & new_nl_ & new_nk_ & new_n_n41_ & new_n_n35_;
  assign new_n_n6_ = ~new_ni0_;
  assign new_nb1_ = new_nc11_ | new_nk12_ | new_nw10_ | new_ns11_ | new_nt11_ | new_ns6_ | new_nk6_ | new_ni2_ | new_nk10_ | new_na9_ | new_nc9_ | new_nw8_ | new_ne6_ | new_nz5_ | new_nj8_;
  assign new_nq1_ = new_ne9_ | new_nd11_ | new_ng11_;
  assign new_n_n67_ = new_nd0_ & new_nw_ & new_n_n38_ & new_n_n2_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_n_n40_;
  assign new_n_n56_ = new_n_n38_ & new_nd0_ & new_na0_ & new_n_n29_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_n_n39_;
  assign new_nx6_ = new_ne0_ & new_ns_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nx_;
  assign new_ni7_ = new_n_n38_ & new_nd0_ & new_n_n7_ & new_n_n16_ & new_n_n15_ & new_nj0_ & new_n_n6_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_nx7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_np0_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_ni8_ = new_nd0_ & new_nc0_ & new_ne0_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_n_n30_;
  assign new_np8_ = new_nc0_ & new_nv_ & new_n_n22_ & new_ns_ & new_nq_ & new_n_n35_ & new_nu_;
  assign new_na9_ = new_nv_ & new_nu_ & new_n_n37_ & new_nz_ & new_ne0_ & new_na_ & new_n_n26_ & new_nk_ & new_n_n41_ & new_n_n35_;
  assign new_n_n7_ = ~new_ng0_;
  assign new_na1_ = new_nb9_ | new_nz10_ | new_np6_ | new_ne6_ | new_nw10_ | new_na9_;
  assign new_na2_ = new_ni8_ | new_no8_ | new_nk8_ | new_ng8_ | new_nf8_;
  assign new_n_n66_ = new_ne0_ & new_n_n37_ & new_n_n29_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_nw_;
  assign new_n_n57_ = new_ne0_ & new_n_n37_ & new_na0_ & new_n_n29_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nc0_;
  assign new_ny6_ = new_ne0_ & new_ns_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nw_;
  assign new_nh7_ = new_n_n38_ & new_nd0_ & new_n_n7_ & new_n_n16_ & new_n_n15_ & new_n_n5_ & new_n_n6_ & new_nk0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_ny7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_nm0_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nh8_ = new_n_n37_ & new_nb0_ & new_n_n38_ & new_n_n32_ & new_nt_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_nq8_ = new_nd0_ & new_n_n39_ & new_n_n38_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_n_n30_;
  assign new_nz8_ = new_nz_ & new_n_n28_ & new_n_n35_ & new_n_n41_ & new_nu_ & new_nv_;
  assign new_n_n8_ = ~new_ns0_;
  assign new_nw0_ = new_nn9_ | new_nm9_;
  assign new_nk1_ = new_ne8_ | new_np9_ | new_ni8_ | new_nf8_ | new_nj9_ | new_no9_ | new_nf9_ | new_ni9_ | new_nq8_ | new_nh7_ | new_ns9_ | new_ng7_ | new_no7_ | new_nx10_ | new_nr9_ | new_ny5_ | new_nm10_ | new_nn7_ | new_nd6_ | new_no12_ | new_nb10_ | new_nr7_ | new_nf6_ | new_nr11_ | new_nx9_ | new_np7_ | new_nc6_ | new_nb11_ | new_nz9_ | new_no11_ | new_ny11_ | new_ng6_ | new_ny9_ | new_nc8_ | new_nu11_ | new_ne11_ | new_nj6_ | new_ny6_ | new_nt6_ | new_ns7_ | new_nd7_ | new_ny10_ | new_nl10_ | new_nw6_ | new_nl9_ | new_ng12_ | new_nm12_ | new_no6_ | new_nx6_ | new_nz11_ | new_na11_ | new_nt9_ | new_nj10_ | new_nr6_ | new_nl12_ | new_nh11_ | new_nh10_ | new_nn1_ | new_nu12_ | new_nx8_ | new_nr8_ | new_nu8_ | new_ny8_ | new_ne9_ | new_no1_ | new_np12_ | new_ni11_ | new_ng10_;
  assign new_nv1_ = new_nr9_ | new_ns9_ | new_nv9_ | new_na7_ | new_nt6_ | new_ni11_ | new_nj10_ | new_nk9_ | new_nz6_ | new_nl9_ | new_np7_ | new_nb10_ | new_nr10_ | new_ns7_ | new_nt9_ | new_nx5_ | new_nb7_ | new_ng7_ | new_nf7_ | new_nm11_ | new_ns10_ | new_nz8_ | new_nj9_ | new_nq9_ | new_ni7_ | new_nf9_ | new_ny8_ | new_nd5_ | new_nu10_ | new_nh7_ | new_na12_ | new_ne7_ | new_np10_ | new_nl7_ | new_nk11_ | new_nh11_ | new_nm7_ | new_nj7_ | new_nb12_ | new_nb11_ | new_nk7_ | new_nq10_;
  assign new_nf2_ = new_n_n49_ | new_n_n48_ | new_n_n59_ | new_n_n43_ | new_n_n52_ | new_n_n54_ | new_n_n53_ | new_n_n68_ | new_n_n67_ | new_ne10_ | new_nl11_ | new_ng9_ | new_n_n44_ | new_n_n55_ | new_n_n45_ | new_n_n65_ | new_n_n63_ | new_n_n66_ | new_n_n62_ | new_n_n64_ | new_n_n51_ | new_n_n60_ | new_n_n61_ | new_n_n56_ | new_n_n50_ | new_n_n57_ | new_n_n47_ | new_n_n58_ | new_n_n46_;
  assign new_n_n58_ = new_nd0_ & new_nc0_ & new_n_n29_ & new_n_n38_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_n_n44_ = new_ne0_ & new_n_n37_ & new_n_n32_ & new_n_n29_ & new_n_n33_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_n_n40_ & new_nc0_;
  assign new_nc6_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_na0_;
  assign new_nn6_ = new_ne0_ & new_n_n37_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_nd7_ = new_ne0_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_n_n39_;
  assign new_no7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_n_n10_ & new_n_n14_ & new_n_n8_ & new_nr0_ & new_n_n11_ & new_n_n12_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nr7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_no0_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nc8_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_nh0_ & new_nj_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nn8_ = new_n_n30_ & new_n_n40_ & new_nd0_ & new_n_n39_ & new_ne0_ & new_na_ & new_ns_ & new_n_n42_ & new_nt_ & new_nu_;
  assign new_ny8_ = new_ne0_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_n_n21_;
  assign new_nx9_ = new_n_n38_ & new_ns_ & new_nu_ & new_nt_ & new_nv_ & new_nd0_;
  assign new_ni10_ = new_n_n38_ & new_n_n37_ & new_ns_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nc0_;
  assign new_n_n1_ = ~new_nm_;
  assign new_ng1_ = new_ni8_ | new_nw6_ | new_nv10_ | new_ne12_ | new_nv6_ | new_nr11_ | new_nh8_ | new_nh6_ | new_no11_ | new_nz7_ | new_nj6_ | new_nu8_ | new_np9_ | new_na11_ | new_nw7_ | new_no9_ | new_nr8_ | new_no1_ | new_no12_ | new_nv7_ | new_nn6_ | new_ns12_ | new_ng6_ | new_nu7_ | new_nt7_ | new_nr6_ | new_np12_ | new_ny5_ | new_nj12_ | new_nq7_ | new_nn1_ | new_ni12_ | new_nd6_ | new_nl9_ | new_nt9_ | new_np11_ | new_nc12_ | new_nb10_ | new_ny6_ | new_nn12_ | new_nm12_ | new_nc6_ | new_nx6_;
  assign new_nl1_ = new_np9_ | new_no6_ | new_nf10_ | new_ng10_ | new_ny9_ | new_nl10_ | new_nj10_ | new_nl12_ | new_nm12_ | new_nj7_ | new_nv6_ | new_ni7_ | new_ny6_ | new_nu11_ | new_nn6_ | new_ni12_ | new_nh7_ | new_nj12_ | new_np11_ | new_ng12_ | new_nx9_ | new_ng7_ | new_nf6_ | new_nn12_ | new_nx10_ | new_nh6_ | new_nv10_ | new_nc12_ | new_ne12_ | new_nb7_ | new_nd7_ | new_nh8_ | new_nu12_ | new_nu8_ | new_ni9_ | new_no9_ | new_nf8_ | new_nx8_ | new_nr8_ | new_np12_ | new_nz11_ | new_ne8_ | new_ns12_ | new_ny11_;
  assign new_nu1_ = new_nd10_ | new_nq11_ | new_nf12_ | new_ng8_ | new_nx11_ | new_nc10_ | new_nk12_ | new_nt12_ | new_no8_ | new_nk8_ | new_nu9_;
  assign new_n_n68_ = new_n_n29_ & new_ne0_ & new_n_n41_ & new_nv_ & new_nt_ & new_nc0_ & new_n_n37_;
  assign new_n_n59_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_n_n2_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_n_n54_ = new_n_n38_ & new_nd0_ & new_nx_ & new_n_n29_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_n_n39_;
  assign new_nd6_ = new_n_n37_ & new_nc0_ & new_n_n38_ & new_ns_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_na0_;
  assign new_nm6_ = new_ne0_ & new_n_n37_ & new_na_ & new_nt_ & new_n_n41_ & new_nv_ & new_nc0_;
  assign new_ne7_ = new_nc0_ & new_nv_ & new_ni_ & new_ns_ & new_nq_ & new_n_n35_ & new_nu_;
  assign new_nn7_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_ns7_ = new_ne0_ & new_nc0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nw_;
  assign new_nb8_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_nf0_ & new_nj_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_no8_ = new_n_n39_ & new_n_n30_ & new_ne0_ & new_nd0_ & new_nf_ & new_nt_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_nx8_ = new_n_n38_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_n_n21_;
  assign new_ny9_ = new_nd0_ & new_n_n39_ & new_n_n38_ & new_n_n41_ & new_nu_ & new_nt_ & new_nv_ & new_nw_;
  assign new_nh10_ = new_ne0_ & new_nd0_ & new_ns_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_n_n39_;
  assign new_n_n2_ = ~new_nb_;
  assign new_nt0_ = new_nl6_ | new_nn9_ | new_ne10_ | new_nl11_ | new_nm9_ | new_ng9_;
  assign new_nf1_ = new_ns9_ | new_nz9_ | new_nt6_ | new_nr9_ | new_no6_ | new_nj9_ | new_nj6_ | new_nl12_ | new_ng6_ | new_nd7_ | new_nd11_ | new_ne11_ | new_ny9_ | new_nm10_ | new_ni12_ | new_nl9_ | new_nf6_ | new_nl10_ | new_np7_ | new_nh10_ | new_nq7_ | new_nr11_ | new_ng11_ | new_nt9_ | new_nd6_ | new_nn12_ | new_nn1_ | new_nx8_ | new_nd8_ | new_nf9_ | new_ni9_ | new_ny8_ | new_ne9_ | new_ny10_ | new_no1_ | new_nx9_ | new_nf8_ | new_nb10_ | new_nx10_ | new_ny5_ | new_nh11_ | new_ng10_ | new_nu12_ | new_nb11_ | new_nm8_ | new_nu11_ | new_ni8_ | new_nr6_ | new_ny11_ | new_na11_ | new_nh8_ | new_ng12_;
  assign new_nm1_ = new_ny9_ | new_ng10_ | new_no6_ | new_nf10_ | new_nd11_ | new_nl10_ | new_nd7_ | new_nl12_ | new_nx10_ | new_nw6_ | new_nx6_ | new_ne12_ | new_nm8_ | new_ni12_ | new_nu11_ | new_ng12_ | new_np11_ | new_nh8_ | new_nj12_ | new_nf8_ | new_nv6_ | new_ne8_ | new_nn6_ | new_nm12_ | new_nx9_ | new_ns7_ | new_no12_ | new_nc12_ | new_ng11_ | new_nr6_ | new_nv10_ | new_nc6_ | new_na12_ | new_no7_ | new_no11_ | new_nl7_ | new_nh6_ | new_nf6_ | new_nx8_ | new_ni7_ | new_no9_ | new_np9_ | new_ne9_ | new_ni9_ | new_nd5_ | new_nd6_ | new_np12_ | new_nk7_ | new_nu12_ | new_ny11_;
  assign new_nx1_ = new_nq12_ | new_np6_ | new_ne6_ | new_nj8_ | new_nk6_ | new_ns11_;
  assign new_ne2_ = new_nl8_ | new_nx8_ | new_nc8_ | new_nk7_ | new_nt7_ | new_nw8_ | new_nb8_ | new_nm8_ | new_nu7_ | new_nz8_ | new_nj7_ | new_nb6_ | new_nn6_ | new_nv7_ | new_ny8_ | new_nm7_ | new_no1_ | new_nw7_ | new_nf6_ | new_nl7_ | new_ng6_ | new_ns6_ | new_ng8_ | new_nq8_ | new_na9_ | new_nc6_ | new_nq6_ | new_ne12_ | new_nn1_ | new_nf8_ | new_np6_ | new_ne8_ | new_nn8_ | new_nr7_ | new_nr6_ | new_ni7_ | new_ne6_ | new_nd8_ | new_no8_ | new_ns7_ | new_na11_ | new_nh7_ | new_nl9_ | new_na12_ | new_nd10_ | new_nq12_ | new_nf12_ | new_ni6_ | new_nk8_ | new_na6_ | new_nz10_ | new_nc10_ | new_nt9_ | new_nb12_ | new_ng12_ | new_nq11_ | new_nh6_ | new_nj8_ | new_nd6_ | new_ny10_ | new_nu11_ | new_nh11_ | new_nc12_ | new_nu6_ | new_nn11_ | new_nk6_ | new_ni8_ | new_ny5_ | new_ni11_ | new_nx10_ | new_nt11_ | new_nh12_ | new_nd12_ | new_nv6_ | new_nz5_ | new_nj6_ | new_nh8_ | new_nn9_ | new_nc9_ | new_nw10_ | new_nx9_ | new_nf11_ | new_nx11_ | new_nx7_ | new_nn12_ | new_no7_ | new_nb9_ | new_nf7_ | new_no9_ | new_ng11_ | new_np8_ | new_nk11_ | new_nm10_ | new_nw11_ | new_nt6_ | new_nm9_ | new_nk9_ | new_nj11_ | new_nn10_ | new_ni12_ | new_nl6_ | new_ns11_ | new_nv9_ | new_no10_ | new_nc7_ | new_nd7_ | new_nr11_ | new_nv10_ | new_nj9_ | new_ng10_ | new_nm6_ | new_np10_ | new_no11_ | new_np12_ | new_no6_ | new_ni9_ | new_nf10_ | new_nj12_ | new_nx5_ | new_ns12_ | new_nr8_ | new_nb7_ | new_nu9_ | new_nq10_ | new_nt12_ | new_nu12_ | new_nv12_ | new_nz6_ | new_ny6_ | new_no12_ | new_nt8_ | new_nw6_ | new_nv8_ | new_nz1_ | new_nx6_ | new_nr12_ | new_ns8_ | new_ny11_ | new_nt10_ | new_nm12_ | new_nn7_ | new_ny7_ | new_ng7_ | new_nh10_ | new_ni2_ | new_nu10_ | new_np11_ | new_nd11_ | new_nd5_ | new_nz7_ | new_nl12_ | new_nq7_ | new_ni10_ | new_nw9_ | new_ne7_ | new_nb10_ | new_ne11_ | new_nz11_ | new_na8_ | new_nk12_ | new_n_n69_ | new_np7_ | new_nh9_ | new_nz9_ | new_nr9_ | new_nj10_ | new_nb11_ | new_ns10_ | new_nf9_ | new_ny9_ | new_ns9_ | new_nd9_ | new_na10_ | new_nq9_ | new_nl10_ | new_nv11_ | new_nm11_ | new_nk10_ | new_nc11_ | new_nr10_ | new_ne9_ | new_na7_ | new_np9_;
  assign new_n_n60_ = new_n_n38_ & new_nd0_ & new_nx_ & new_n_n2_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_n_n40_;
  assign new_n_n53_ = new_ne0_ & new_n_n37_ & new_na0_ & new_n_n29_ & new_nl_ & new_ns_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nc0_;
  assign new_ng2_ = new_ny9_ | new_nl10_ | new_no6_ | new_nx10_ | new_ng10_ | new_nu9_ | new_nd11_ | new_na11_ | new_nd7_ | new_nn1_ | new_ny11_ | new_ng6_ | new_nx9_ | new_ny5_ | new_no1_ | new_nj6_ | new_ng11_ | new_ni12_ | new_nt12_ | new_nk8_ | new_nn12_ | new_nl12_ | new_nx8_ | new_nf8_ | new_no9_ | new_np9_ | new_ne9_ | new_ni9_;
  assign new_nl6_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_nv_ & new_nt_ & new_ny_ & new_n_n39_;
  assign new_nb7_ = new_ne0_ & new_nz_ & new_nk_ & new_n_n35_ & new_ns_ & new_n_n34_ & new_n_n40_;
  assign new_nm7_ = new_n_n38_ & new_nd0_ & new_nf0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_nt7_ = new_nd0_ & new_n_n39_ & new_ne0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nw_;
  assign new_ne8_ = new_nd0_ & new_n_n39_ & new_n_n38_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_nb0_;
  assign new_nl8_ = new_n_n37_ & new_nc0_ & new_ne0_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_n_n30_;
  assign new_nw8_ = new_n_n37_ & new_nw_ & new_ne0_ & new_na_ & new_n_n35_ & new_n_n41_ & new_nu_ & new_nv_;
  assign new_nd9_ = new_na0_ & new_nv_ & new_ne0_ & new_n_n37_ & new_na_ & new_n_n41_ & new_nl_ & new_n_n35_ & new_nu_;
  assign new_no9_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_nb_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_n_n3_ = ~new_nl0_;
  assign new_nu0_ = new_nl11_ | new_ng9_;
  assign new_ne1_ = new_nj9_ | new_no9_ | new_np9_ | new_nr9_ | new_nt6_ | new_ns9_ | new_nb11_ | new_nd11_ | new_no6_ | new_nu12_ | new_ng12_ | new_nh10_ | new_nf6_ | new_nh11_ | new_nx9_ | new_ng10_ | new_nr6_ | new_ne11_ | new_nz9_ | new_nu11_ | new_nm10_ | new_nl10_ | new_no7_ | new_ny11_ | new_ne9_ | new_nx8_ | new_ny8_ | new_nf9_ | new_ni9_ | new_nf8_ | new_nd7_ | new_nx10_ | new_nh8_ | new_nl12_ | new_ny9_ | new_nm8_ | new_ng11_ | new_ny10_ | new_nd6_;
  assign new_nn1_ = new_n_n39_ & new_na0_ & new_ne0_ & new_nd0_ & new_n_n36_ & new_n_n35_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_nw1_ = new_nn8_ | new_ng8_ | new_nc11_ | new_nv12_ | new_nd12_ | new_nk12_ | new_na9_ | new_nc9_ | new_nd9_ | new_nx11_ | new_nb9_ | new_nw8_ | new_nt11_ | new_nf11_ | new_nt10_ | new_nu6_ | new_nb6_ | new_nw10_ | new_ni2_ | new_nz10_ | new_nk10_ | new_nm6_ | new_nf10_ | new_nh9_;
  assign new_n_n69_ = new_ne0_ & new_ns_ & new_nu_ & new_nt_ & new_nv_ & new_na0_;
  assign new_n_n61_ = new_nd_ & new_n_n29_ & new_nb0_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_n_n37_;
  assign new_n_n52_ = new_n_n38_ & new_nd0_ & new_na0_ & new_n_n29_ & new_nr_ & new_ns_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_n_n39_;
  assign new_n_n43_ = new_n_n37_ & new_n_n39_ & new_n_n29_ & new_ne0_ & new_n_n42_ & new_n_n27_ & new_n_n41_ & new_nu_ & new_nt_ & new_nv_ & new_nw_;
  assign new_nb6_ = new_n_n39_ & new_na0_ & new_n_n38_ & new_nd0_ & new_na_ & new_nt_ & new_ns_ & new_n_n34_ & new_n_n40_;
  assign new_nc7_ = new_nw_ & new_nv_ & new_n_n37_ & new_nc0_ & new_n_n38_ & new_n_n23_ & new_n_n41_ & new_n_n25_ & new_nt_ & new_nu_;
  assign new_nl7_ = new_n_n38_ & new_nd0_ & new_ng0_ & new_n_n16_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_nv_ & new_nx_;
  assign new_nu7_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_n_n13_ & new_n_n12_ & new_nn0_ & new_nq0_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nd8_ = new_n_n39_ & new_nw_ & new_ne0_ & new_n_n37_ & new_n_n17_ & new_n_n35_ & new_n_n41_ & new_n_n34_ & new_nv_;
  assign new_nm8_ = new_n_n37_ & new_nc0_ & new_n_n38_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_n_n30_;
  assign new_nv8_ = new_n_n38_ & new_n_n37_ & new_nn_ & new_n_n40_ & new_n_n20_ & new_n_n30_ & new_n_n39_;
  assign new_ne9_ = new_n_n38_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_nv_ & new_na0_;
  assign new_nn9_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_nv_ & new_nt_ & new_na0_ & new_n_n39_;
  assign new_n_n4_ = ~new_nk0_;
  assign new_nw10_ = new_n_n35_ & new_ns_ & new_nv_ & new_nu_ & new_nz_ & new_n_n37_ & new_n_n39_ & new_ne0_ & new_na_ & new_nk_ & new_n_n42_ & new_n_n26_ & new_n_n27_;
  assign new_nh11_ = new_n_n39_ & new_na0_ & new_ne0_ & new_nd0_ & new_nl_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_ns11_ = new_nc0_ & new_nw_ & new_n_n38_ & new_nd0_ & new_na_ & new_nt_ & new_n_n41_ & new_nu_ & new_n_n40_;
  assign new_nd12_ = new_n_n39_ & new_nx_ & new_n_n38_ & new_nd0_ & new_na_ & new_n_n35_ & new_n_n41_ & new_nu_ & new_n_n40_;
  assign new_no12_ = new_nc0_ & new_nw_ & new_ne0_ & new_n_n37_ & new_nd_ & new_nt_ & new_n_n41_ & new_nu_ & new_n_n40_;
  assign new_nv10_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nx_;
  assign new_ni11_ = new_ne0_ & new_ns_ & new_n_n34_ & new_nt_ & new_nv_ & new_nw_;
  assign new_nr11_ = new_nd0_ & new_nc0_ & new_ne0_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_ne12_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_ns_ & new_nu_ & new_nt_ & new_n_n40_ & new_n_n30_;
  assign new_nn12_ = new_nd0_ & new_nw_ & new_n_n38_ & new_nb_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_n_n40_;
  assign new_nu10_ = new_nc0_ & new_nv_ & new_nh_ & new_ns_ & new_n_n25_ & new_n_n35_ & new_nu_;
  assign new_nj11_ = new_n_n38_ & new_n_n37_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nc0_;
  assign new_nu11_ = new_ne0_ & new_nd0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_n_n40_ & new_n_n39_;
  assign new_nb12_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_na0_;
  assign new_nm12_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_n_n34_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_nt10_ = new_ne0_ & new_n_n37_ & new_na_ & new_nt_ & new_ns_ & new_nu_ & new_nv_;
  assign new_nk11_ = new_ne0_ & new_nz_ & new_n_n28_ & new_nt_ & new_ns_ & new_n_n34_ & new_nv_;
  assign new_nt11_ = new_n_n40_ & new_n_n34_ & new_nd0_ & new_n_n39_ & new_n_n38_ & new_na_ & new_n_n42_ & new_n_n32_ & new_n_n41_ & new_n_n35_;
  assign new_nc12_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nx_;
  assign new_nl12_ = new_n_n38_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_nc0_;
  assign new_n_n0_ = ~new_nn_;
  assign new_ns10_ = new_nu_ & new_n_n35_ & new_nz_ & new_nv_ & new_n_n39_ & new_ne0_ & new_n_n37_ & new_na_ & new_n_n28_ & new_n_n42_ & new_n_n27_ & new_ns_;
  assign new_nv12_ = new_nw_ & new_n_n40_ & new_nd0_ & new_n_n39_ & new_n_n38_ & new_na_ & new_n_n41_ & new_n_n42_ & new_nt_ & new_nu_;
  assign new_n_n32_ = ~new_nd_;
  assign new_n_n21_ = ~new_na0_;
  assign new_n_n10_ = ~new_no0_;
  assign new_nr10_ = new_nz_ & new_nv_ & new_n_n37_ & new_n_n39_ & new_ne0_ & new_nf_ & new_ns_ & new_n_n28_ & new_n_n35_ & new_nu_;
  assign new_n_n42_ = ~new_nf_;
  assign new_n_n33_ = ~new_nc_;
  assign new_n_n20_ = ~new_no_;
  assign new_n_n11_ = ~new_nq0_;
  assign new_n_n41_ = ~new_ns_;
  assign new_n_n30_ = ~new_nb0_;
  assign new_n_n23_ = ~new_nh_;
  assign new_n_n12_ = ~new_np0_;
  assign new_n_n40_ = ~new_nv_;
  assign new_n_n31_ = ~new_ng_;
  assign new_n_n22_ = ~new_ni_;
  assign new_n_n13_ = ~new_nm0_;
  assign new_nv11_ = new_n_n38_ & new_n_n37_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_n_n40_ & new_nc0_;
  assign new_ng12_ = new_n_n39_ & new_na0_ & new_n_n38_ & new_nd0_ & new_nr_ & new_n_n35_ & new_ns_ & new_nu_ & new_n_n40_;
  assign new_nr12_ = new_n_n37_ & new_nc0_ & new_n_n38_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_n_n36_ = ~new_nr_;
  assign new_n_n25_ = ~new_nq_;
  assign new_n_n14_ = ~new_nn0_;
  assign new_nw11_ = new_nc0_ & new_n_n40_ & new_ne0_ & new_n_n37_ & new_n_n33_ & new_n_n41_ & new_n_n32_ & new_n_n35_ & new_n_n34_;
  assign new_nf12_ = new_n_n40_ & new_nu_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_n_n33_ & new_ng_ & new_n_n32_ & new_n_n41_ & new_n_n35_;
  assign new_ns12_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_na0_;
  assign new_n_n37_ = ~new_nd0_;
  assign new_n_n24_ = ~new_nz_;
  assign new_n_n15_ = ~new_nh0_;
  assign new_nb11_ = new_n_n39_ & new_nz_ & new_ne0_ & new_nd0_ & new_nl_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_nm11_ = new_ne0_ & new_ns_ & new_nu_ & new_nt_ & new_nv_ & new_nw_;
  assign new_nt12_ = new_n_n39_ & new_nw_ & new_n_n38_ & new_nd0_ & new_nf_ & new_nt_ & new_n_n41_ & new_nu_ & new_n_n40_;
  assign new_n_n34_ = ~new_nu_;
  assign new_n_n27_ = ~new_np_;
  assign new_n_n16_ = ~new_nf0_;
  assign new_nc11_ = new_nu_ & new_n_n35_ & new_na0_ & new_nv_ & new_n_n39_ & new_ne0_ & new_n_n37_ & new_na_ & new_n_n26_ & new_n_n42_ & new_n_n27_ & new_ns_;
  assign new_nl11_ = new_n_n37_ & new_ny_ & new_ne0_ & new_n_n29_ & new_nt_ & new_ns_ & new_nu_ & new_nv_;
  assign new_nu12_ = new_nd0_ & new_n_n39_ & new_ne0_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_n_n35_ = ~new_nt_;
  assign new_n_n26_ = ~new_nl_;
  assign new_n_n17_ = ~new_nj_;
  assign new_na11_ = new_n_n39_ & new_nz_ & new_n_n38_ & new_nd0_ & new_nl_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_nd11_ = new_n_n39_ & new_na0_ & new_n_n38_ & new_nd0_ & new_n_n26_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_no11_ = new_nw_ & new_n_n40_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_n_n33_ & new_n_n41_ & new_n_n32_ & new_nt_ & new_nu_;
  assign new_nz11_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_ny_;
  assign new_nk12_ = new_n_n40_ & new_nu_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_na_ & new_n_n32_ & new_n_n33_ & new_n_n41_ & new_n_n35_;
  assign new_n_n29_ = ~new_na_;
  assign new_n_n18_ = ~new_ne_;
  assign new_nz10_ = new_n_n35_ & new_ns_ & new_nv_ & new_nu_ & new_nz_ & new_n_n37_ & new_n_n39_ & new_ne0_ & new_na_ & new_nk_ & new_n_n42_ & new_nl_ & new_n_n27_;
  assign new_ne11_ = new_n_n39_ & new_na0_ & new_ne0_ & new_nd0_ & new_n_n26_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_nn11_ = new_n_n40_ & new_nu_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n41_ & new_n_n35_;
  assign new_na12_ = new_n_n38_ & new_nd0_ & new_n_n41_ & new_nu_ & new_n_n35_ & new_n_n40_ & new_ny_;
  assign new_nj12_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_nw_;
  assign new_n_n28_ = ~new_nk_;
  assign new_n_n19_ = ~new_nx_;
  assign new_ny10_ = new_n_n39_ & new_nz_ & new_ne0_ & new_nd0_ & new_n_n26_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_nf11_ = new_nu_ & new_n_n35_ & new_na0_ & new_nv_ & new_n_n39_ & new_ne0_ & new_n_n37_ & new_na_ & new_nl_ & new_n_n42_ & new_n_n27_ & new_ns_;
  assign new_nq11_ = new_nc0_ & new_n_n40_ & new_ne0_ & new_n_n37_ & new_nd_ & new_n_n41_ & new_ng_ & new_n_n35_ & new_nu_;
  assign new_nx11_ = new_n_n40_ & new_n_n34_ & new_n_n37_ & new_nc0_ & new_ne0_ & new_na_ & new_n_n32_ & new_nc_ & new_n_n41_ & new_n_n35_;
  assign new_ni12_ = new_nd0_ & new_nx_ & new_n_n38_ & new_nb_ & new_nt_ & new_n_n41_ & new_n_n34_ & new_n_n40_;
  assign new_np12_ = new_n_n37_ & new_n_n39_ & new_ne0_ & new_n_n41_ & new_nu_ & new_nt_ & new_n_n40_ & new_nx_;
  assign new_n_n38_ = ~new_ne0_;
  assign new_nx10_ = new_n_n39_ & new_nz_ & new_n_n38_ & new_nd0_ & new_n_n26_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_ng11_ = new_n_n39_ & new_na0_ & new_n_n38_ & new_nd0_ & new_nl_ & new_n_n35_ & new_ns_ & new_nu_ & new_nv_;
  assign new_np11_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_n_n40_ & new_n_n39_;
  assign new_ny11_ = new_n_n38_ & new_nd0_ & new_n_n41_ & new_n_n34_ & new_n_n35_ & new_n_n40_ & new_nc0_;
  assign new_nh12_ = new_nc0_ & new_n_n40_ & new_ne0_ & new_n_n37_ & new_nd_ & new_n_n41_ & new_n_n31_ & new_n_n35_ & new_nu_;
  assign new_nq12_ = new_na0_ & new_n_n40_ & new_nd0_ & new_n_n39_ & new_n_n38_ & new_na_ & new_ns_ & new_n_n36_ & new_n_n35_ & new_nu_;
  assign new_n_n39_ = ~new_nc0_;
endmodule


