// Benchmark "top" written by ABC on Fri Mar 31 12:10:25 2023

module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0,
    pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0, pb, pr0, pc,
    ps0, pd, pt0, pe, pu0, pf, pv0, pg, pw0, ph, px0, pi, py0, pj, pz0, pk,
    pl, pm, pn, po,
    pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pg2, pd2, pg1, pe2, pf1,
    pi1, ph1, ph2, pk1, pi2, pj1, pm1, pl1, po1, pn1, pq1, pp1, ps1, pr1,
    pu1, pt1, pw1, pv1, py1, px1, pz1  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0,
    pw, ph0, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0, pb,
    pr0, pc, ps0, pd, pt0, pe, pu0, pf, pv0, pg, pw0, ph, px0, pi, py0, pj,
    pz0, pk, pl, pm, pn, po;
  output pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pg2, pd2, pg1, pe2, pf1,
    pi1, ph1, ph2, pk1, pi2, pj1, pm1, pl1, po1, pn1, pq1, pp1, ps1, pr1,
    pu1, pt1, pw1, pv1, py1, px1, pz1;
  wire new_np_, new_na0_, new_nq_, new_nb0_, new_nr_, new_nc0_, new_ns_,
    new_nd0_, new_nt_, new_ne0_, new_nu_, new_nf0_, new_nv_, new_ng0_,
    new_nw_, new_nh0_, new_ni0_, new_ny_, new_nj0_, new_nz_, new_nk0_,
    new_nl0_, new_nm0_, new_nn0_, new_no0_, new_np0_, new_na_, new_nq0_,
    new_nb_, new_nr0_, new_nc_, new_ns0_, new_nd_, new_nt0_, new_ne_,
    new_nu0_, new_nf_, new_nv0_, new_ng_, new_nw0_, new_nh_, new_nx0_,
    new_ni_, new_ny0_, new_nj_, new_nz0_, new_nk_, new_nl_, new_nm_,
    new_nn_, new_no_, new_n_n330_, new_n_n322_, new_n_n313_, new_n_n303_,
    new_n_n292_, new_n_n281_, new_nl1_, new_n_n240_, new_nm1_, new_n_n220_,
    new_n_n211_, new_n_n202_, new_n_n196_, new_n_n155_, new_n_n146_,
    new_n_n136_, new_n_n125_, new_n_n114_, new_n_n103_, new_nb1_, new_nd1_,
    new_n_n312_, new_n_n304_, new_n_n291_, new_n_n282_, new_n_n260_,
    new_n_n239_, new_n_n230_, new_no1_, new_n_n212_, new_nx1_, new_nb2_,
    new_n_n154_, new_ns1_, new_n_n135_, new_n_n126_, new_n_n113_,
    new_n_n104_, new_n_n332_, new_n_n323_, new_n_n311_, new_n_n301_,
    new_n_n294_, new_n_n283_, new_n_n259_, new_n_n249_, new_n_n231_,
    new_n_n219_, new_n_n209_, new_nw1_, new_na2_, new_n_n175_, new_n_n164_,
    new_n_n134_, new_n_n123_, new_n_n116_, new_n_n105_, new_n_n331_,
    new_n_n324_, new_n_n310_, new_n_n302_, new_n_n293_, new_n_n284_,
    new_n_n258_, new_n_n250_, new_n_n241_, new_n_n218_, new_n_n210_,
    new_n_n203_, new_nz1_, new_n_n174_, new_n_n165_, new_n_n133_,
    new_n_n124_, new_n_n115_, new_n_n106_, new_n_n309_, new_n_n299_,
    new_n_n278_, new_n_n268_, new_n_n217_, new_nv1_, new_n_n199_, new_nd2_,
    new_n_n183_, new_n_n132_, new_n_n121_, new_n_n110_, new_n_n99_,
    new_n_n9_, new_ng1_, new_n_n300_, new_n_n277_, new_n_n269_,
    new_n_n216_, new_n_n208_, new_n_n193_, new_n_n192_, new_n_n184_,
    new_n_n131_, new_n_n122_, new_n_n109_, new_n_n100_, new_n_n290_,
    new_nh1_, new_n_n270_, new_n_n215_, new_n_n201_, new_n_n194_,
    new_n_n130_, new_n_n119_, new_n_n112_, new_n_n101_, new_n_n289_,
    new_n_n280_, new_n_n279_, new_n_n207_, new_n_n200_, new_n_n195_,
    new_n_n129_, new_n_n120_, new_n_n111_, new_n_n102_, new_n_n333_,
    new_n_n275_, new_n_n264_, new_n_n253_, new_n_n243_, new_n_n232_,
    new_n_n189_, new_n_n179_, new_n_n169_, new_n_n158_, new_n_n148_,
    new_n_n139_, new_n_n5_, new_n_n334_, new_n_n274_, new_n_n265_,
    new_n_n252_, new_n_n244_, new_n_n224_, new_n_n188_, new_n_n180_,
    new_n_n168_, new_n_n159_, new_n_n147_, new_n_n140_, new_n_n6_,
    new_n_n325_, new_n_n317_, new_n_n276_, new_n_n266_, new_n_n251_,
    new_n_n234_, new_n_n225_, new_n_n191_, new_n_n181_, new_n_n167_,
    new_n_n156_, new_n_n150_, new_n_n141_, new_n_n7_, new_nc1_,
    new_n_n318_, new_nk1_, new_n_n267_, new_n_n242_, new_n_n233_,
    new_n_n226_, new_n_n190_, new_n_n182_, new_n_n166_, new_n_n157_,
    new_n_n149_, new_nh2_, new_n_n8_, new_na1_, new_n_n327_, new_ne1_,
    new_n_n316_, new_n_n307_, new_n_n296_, new_n_n285_, new_n_n271_,
    new_n_n257_, new_n_n247_, new_n_n236_, new_n_n227_, new_n_n214_,
    new_n_n205_, new_n_n197_, new_ne2_, new_n_n176_, new_n_n173_,
    new_n_n162_, new_n_n151_, new_n_n142_, new_n_n118_, new_n_n107_,
    new_n_n1_, new_n_n326_, new_n_n319_, new_n_n315_, new_n_n308_,
    new_n_n295_, new_n_n286_, new_n_n261_, new_n_n256_, new_n_n248_,
    new_n_n235_, new_nn1_, new_n_n223_, new_n_n204_, new_n_n198_,
    new_n_n185_, new_n_n177_, new_n_n172_, new_n_n163_, new_ng2_,
    new_n_n143_, new_n_n117_, new_n_n108_, new_n_n2_, new_n_n335_,
    new_n_n329_, new_n_n320_, new_n_n314_, new_n_n305_, new_n_n298_,
    new_n_n287_, new_n_n273_, new_n_n262_, new_n_n255_, new_n_n245_,
    new_n_n238_, new_n_n228_, new_n_n222_, new_nr1_, new_ny1_, new_n_n187_,
    new_nf2_, new_n_n171_, new_n_n160_, new_n_n153_, new_n_n144_,
    new_n_n138_, new_n_n127_, new_n_n3_, new_n_n336_, new_n_n328_,
    new_n_n321_, new_nf1_, new_n_n306_, new_n_n297_, new_n_n288_,
    new_n_n272_, new_n_n263_, new_n_n254_, new_n_n246_, new_n_n237_,
    new_n_n229_, new_n_n221_, new_n_n213_, new_n_n206_, new_n_n186_,
    new_n_n178_, new_n_n170_, new_n_n161_, new_n_n152_, new_n_n145_,
    new_n_n137_, new_n_n128_, new_n_n4_, new_n_n93_, new_n_n82_,
    new_n_n71_, new_n_n60_, new_ni2_, new_n_n94_, new_n_n81_, new_n_n72_,
    new_n_n59_, new_n_n50_, new_n_n95_, new_n_n80_, new_n_n69_, new_n_n62_,
    new_n_n51_, new_n_n96_, new_n_n79_, new_n_n70_, new_n_n61_, new_n_n52_,
    new_n_n0_, new_n_n97_, new_n_n43_, new_n_n32_, new_n_n21_, new_n_n10_,
    new_n_n98_, new_n_n42_, new_n_n33_, new_n_n20_, new_n_n11_, new_n_n41_,
    new_n_n30_, new_n_n23_, new_n_n12_, new_n_n40_, new_n_n31_, new_n_n22_,
    new_n_n13_, new_n_n68_, new_n_n57_, new_n_n47_, new_n_n36_, new_n_n25_,
    new_n_n14_, new_n_n67_, new_n_n58_, new_n_n46_, new_n_n37_, new_n_n24_,
    new_n_n15_, new_n_n88_, new_n_n77_, new_n_n45_, new_n_n34_, new_n_n27_,
    new_n_n16_, new_n_n87_, new_n_n78_, new_n_n44_, new_n_n35_, new_n_n26_,
    new_n_n17_, new_n_n89_, new_n_n86_, new_n_n75_, new_n_n64_, new_n_n53_,
    new_n_n29_, new_n_n18_, new_n_n90_, new_n_n85_, new_n_n76_, new_n_n63_,
    new_n_n54_, new_n_n28_, new_n_n19_, new_n_n91_, new_n_n84_, new_n_n73_,
    new_n_n66_, new_n_n55_, new_n_n49_, new_n_n38_, new_n_n92_, new_n_n83_,
    new_n_n74_, new_n_n65_, new_n_n56_, new_n_n48_, new_n_n39_;
  assign pa1 = new_na1_;
  assign pb2 = new_nb2_;
  assign new_np_ = pp;
  assign new_na0_ = pa0;
  assign pc2 = new_nh0_;
  assign new_nq_ = pq;
  assign new_nb0_ = pb0;
  assign pc1 = new_nc1_;
  assign new_nr_ = pr;
  assign pa2 = new_na2_;
  assign pb1 = new_nb1_;
  assign new_nc0_ = pc0;
  assign new_ns_ = ps;
  assign new_nd0_ = pd0;
  assign pe1 = new_ne1_;
  assign pf2 = new_nf2_;
  assign new_nt_ = pt;
  assign pd1 = new_nd1_;
  assign new_ne0_ = pe0;
  assign pg2 = new_ng2_;
  assign new_nu_ = pu;
  assign pd2 = new_nd2_;
  assign new_nf0_ = pf0;
  assign pg1 = new_ng1_;
  assign new_nv_ = pv;
  assign pe2 = new_ne2_;
  assign pf1 = new_nf1_;
  assign new_ng0_ = pg0;
  assign new_nw_ = pw;
  assign new_nh0_ = ph0;
  assign pi1 = new_nm0_;
  assign ph1 = new_nh1_;
  assign new_ni0_ = pi0;
  assign new_ny_ = py;
  assign ph2 = new_nh2_;
  assign new_nj0_ = pj0;
  assign pk1 = new_nk1_;
  assign new_nz_ = pz;
  assign pi2 = new_ni2_;
  assign pj1 = new_nn0_;
  assign new_nk0_ = pk0;
  assign new_nl0_ = pl0;
  assign pm1 = new_nm1_;
  assign pl1 = new_nl1_;
  assign new_nm0_ = pm0;
  assign new_nn0_ = pn0;
  assign po1 = new_no1_;
  assign pn1 = new_nn1_;
  assign new_no0_ = po0;
  assign new_np0_ = pp0;
  assign pq1 = new_nz_;
  assign new_na_ = pa;
  assign pp1 = new_ny_;
  assign new_nq0_ = pq0;
  assign new_nb_ = pb;
  assign new_nr0_ = pr0;
  assign ps1 = new_ns1_;
  assign new_nc_ = pc;
  assign pr1 = new_nr1_;
  assign new_ns0_ = ps0;
  assign new_nd_ = pd;
  assign new_nt0_ = pt0;
  assign pu1 = new_ny0_;
  assign new_ne_ = pe;
  assign pt1 = new_nx0_;
  assign new_nu0_ = pu0;
  assign new_nf_ = pf;
  assign new_nv0_ = pv0;
  assign pw1 = new_nw1_;
  assign new_ng_ = pg;
  assign pv1 = new_nv1_;
  assign new_nw0_ = pw0;
  assign new_nh_ = ph;
  assign new_nx0_ = px0;
  assign py1 = new_ny1_;
  assign new_ni_ = pi;
  assign px1 = new_nx1_;
  assign new_ny0_ = py0;
  assign new_nj_ = pj;
  assign new_nz0_ = pz0;
  assign new_nk_ = pk;
  assign pz1 = new_nz1_;
  assign new_nl_ = pl;
  assign new_nm_ = pm;
  assign new_nn_ = pn;
  assign new_no_ = po;
  assign new_n_n330_ = new_n_n38_ & new_n_n24_ & new_na0_ & new_n_n19_;
  assign new_n_n322_ = new_nc0_ & new_nv_;
  assign new_n_n313_ = new_n_n8_ & new_n_n18_ & new_nq0_;
  assign new_n_n303_ = new_n_n26_ & new_np0_ & new_n_n18_ & new_n_n41_ & new_nv_ & new_n_n37_ & new_n_n19_;
  assign new_n_n292_ = new_n_n1_ & new_n_n26_ & new_n_n41_ & new_n_n37_ & new_ng_ & new_n_n6_ & new_np0_;
  assign new_n_n281_ = new_np0_ & new_n_n37_ & new_n_n1_ & new_n_n36_ & new_n_n40_ & new_n_n24_ & new_n_n7_ & new_n_n41_ & new_n_n8_;
  assign new_nl1_ = new_n_n245_ | new_n_n244_ | new_n_n242_ | new_n_n241_ | new_n_n243_ | new_n_n230_ | new_n_n239_ | new_n_n240_ | new_n_n236_ | new_n_n235_ | new_n_n238_ | new_n_n237_ | new_n_n231_ | new_n_n233_ | new_n_n232_ | new_n_n234_ | new_n_n248_ | new_n_n250_ | new_n_n249_ | new_n_n247_ | new_n_n246_;
  assign new_n_n240_ = new_no_ & new_nq_ & new_nq0_ & new_np_;
  assign new_nm1_ = new_n_n228_ | new_n_n229_;
  assign new_n_n220_ = new_n_n3_ & new_n_n4_ & new_nd_ & new_n_n8_ & new_np0_ & new_n_n41_ & new_nc_ & new_n_n24_ & new_n_n40_ & new_n_n5_;
  assign new_n_n211_ = new_n_n41_ & new_n_n26_ & new_ni0_ & new_n_n37_;
  assign new_n_n202_ = new_nr_ & new_ns_ & new_nk0_;
  assign new_n_n196_ = new_n_n24_ & new_n_n4_ & new_ne0_ & new_n_n3_ & new_n_n41_ & new_n_n40_ & new_n_n5_ & new_no_ & new_n_n7_;
  assign new_n_n155_ = new_n_n12_ & new_n_n13_ & new_n_n11_ & new_nd_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_n_n17_ & new_n_n16_ & new_n_n30_ & new_n_n15_ & new_n_n14_;
  assign new_n_n146_ = new_nh_ & new_n_n18_ & new_ne0_;
  assign new_n_n136_ = new_n_n22_ & new_n_n31_ & new_n_n30_ & new_n_n23_ & new_n_n38_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n125_ = new_n_n23_ & new_n_n31_ & new_na_ & new_n_n30_ & new_n_n38_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n114_ = new_n_n25_ & new_n_n31_ & new_nn_ & new_n_n23_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n103_ = new_n_n32_ & new_n_n33_ & new_n_n25_ & new_n_n31_ & new_n_n30_ & new_n_n36_ & new_n_n21_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_nb1_ = new_n_n327_ | new_n_n329_ | new_n_n328_ | new_n_n326_ | new_n_n325_;
  assign new_nd1_ = new_n_n319_ | new_n_n321_ | new_n_n320_ | new_n_n322_;
  assign new_n_n312_ = new_n_n8_ & new_nq0_ & new_n_n6_;
  assign new_n_n304_ = new_ng_ & new_nd0_ & new_n_n40_ & new_np_ & new_no_ & new_nu_ & new_n_n24_;
  assign new_n_n291_ = new_n_n37_ & new_n_n8_ & new_np0_ & new_n_n19_ & new_n_n40_ & new_n_n24_ & new_n_n18_ & new_n_n41_ & new_n_n25_;
  assign new_n_n282_ = new_np0_ & new_n_n37_ & new_n_n1_ & new_n_n36_ & new_n_n40_ & new_n_n24_ & new_n_n18_ & new_n_n41_ & new_n_n8_;
  assign new_n_n260_ = new_nj0_ & new_na_;
  assign new_n_n239_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_nu_ & new_n_n8_ & new_n_n24_;
  assign new_n_n230_ = new_no_ & new_n_n8_ & new_n_n24_ & new_np_ & new_n_n37_ & new_ne_ & new_nd0_ & new_n_n41_ & new_n_n36_;
  assign new_no1_ = new_n_n217_ | new_n_n216_ | new_n_n192_ | new_n_n218_ | new_n_n215_ | new_n_n214_ | new_n_n219_ | new_n_n213_;
  assign new_n_n212_ = new_nj0_ & new_n_n41_;
  assign new_nx1_ = new_n_n201_ | new_nz_ | new_nh0_ | new_n_n200_ | new_n_n199_;
  assign new_nb2_ = new_n_n193_ | new_n_n195_ | new_n_n194_ | new_n_n196_;
  assign new_n_n154_ = new_n_n13_ & new_n_n14_ & new_n_n10_ & new_n_n12_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_no_ & new_n_n17_ & new_n_n23_ & new_n_n16_ & new_n_n15_;
  assign new_ns1_ = new_nh_ & new_nt_ & new_ni0_;
  assign new_n_n135_ = new_n_n25_ & new_n_n31_ & new_n_n30_ & new_n_n23_ & new_n_n21_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n126_ = new_n_n25_ & new_n_n31_ & new_na_ & new_n_n23_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n113_ = new_n_n23_ & new_n_n31_ & new_nn_ & new_n_n30_ & new_n_n38_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n104_ = new_n_n32_ & new_n_n33_ & new_n_n22_ & new_n_n31_ & new_n_n30_ & new_n_n36_ & new_n_n38_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n332_ = new_nf0_ & new_n_n22_;
  assign new_n_n323_ = new_n_n24_ & new_nb0_ & new_n_n40_;
  assign new_n_n311_ = new_n_n18_ & new_nq0_ & new_n_n26_;
  assign new_n_n301_ = new_n_n26_ & new_np0_ & new_n_n18_ & new_ng_ & new_n_n41_ & new_n_n37_ & new_n_n19_;
  assign new_n_n294_ = new_n_n1_ & new_n_n26_ & new_n_n7_ & new_ng_ & new_n_n41_ & new_n_n37_ & new_np0_;
  assign new_n_n283_ = new_n_n6_ & new_n_n37_ & new_n_n1_ & new_np0_ & new_n_n40_ & new_n_n41_ & new_n_n24_ & new_n_n25_ & new_n_n8_;
  assign new_n_n259_ = new_nm_ & new_n_n24_ & new_nd0_;
  assign new_n_n249_ = new_nh0_ & new_ne_;
  assign new_n_n231_ = new_no_ & new_n_n8_ & new_n_n24_ & new_np_ & new_n_n37_ & new_nd0_ & new_nu_ & new_n_n41_ & new_n_n36_;
  assign new_n_n219_ = new_n_n41_ & new_ni_ & new_ni0_ & new_n_n37_;
  assign new_n_n209_ = new_n_n24_ & new_n_n1_ & new_nk0_ & new_n_n41_ & new_n_n38_ & new_nb_ & new_n_n40_ & new_nr_;
  assign new_nw1_ = new_n_n202_ | new_n_n203_;
  assign new_na2_ = new_nr0_ | new_nf0_;
  assign new_n_n175_ = new_n_n15_ & new_n_n16_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_no_ & new_n_n23_ & new_n_n29_ & new_n_n17_ & new_n_n30_;
  assign new_n_n164_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_nb_ & new_nz0_ & new_nl_ & new_n_n23_ & new_n_n30_ & new_n_n17_ & new_n_n16_ & new_n_n15_;
  assign new_n_n134_ = new_n_n25_ & new_n_n22_ & new_n_n30_ & new_n_n23_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n123_ = new_n_n23_ & new_n_n31_ & new_na_ & new_n_n28_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n116_ = new_n_n30_ & new_n_n23_ & new_nm_ & new_n_n28_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n105_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n36_ & new_n_n38_ & new_nh_ & new_n_n21_ & new_n_n35_;
  assign new_n_n331_ = new_nr0_ & new_n_n22_;
  assign new_n_n324_ = new_nb0_ & new_nv_;
  assign new_n_n310_ = new_nq0_ & new_n_n6_ & new_n_n26_;
  assign new_n_n302_ = new_n_n26_ & new_np0_ & new_n_n7_ & new_n_n41_ & new_nv_ & new_n_n37_ & new_n_n19_;
  assign new_n_n293_ = new_n_n1_ & new_n_n26_ & new_nv_ & new_n_n37_ & new_n_n41_ & new_n_n6_ & new_np0_;
  assign new_n_n284_ = new_n_n37_ & new_n_n8_ & new_n_n1_ & new_np0_ & new_n_n40_ & new_n_n24_ & new_n_n7_ & new_n_n41_ & new_n_n25_;
  assign new_n_n258_ = new_nm_ & new_n_n24_ & new_np0_;
  assign new_n_n250_ = new_nh0_ & new_nu_;
  assign new_n_n241_ = new_no_ & new_nq_ & new_np0_ & new_np_;
  assign new_n_n218_ = new_n_n6_ & new_n_n41_ & new_n_n24_ & new_ni_ & new_np0_ & new_ng_;
  assign new_n_n210_ = new_na_ & new_n_n26_ & new_n_n37_ & new_ni0_ & new_n_n10_;
  assign new_n_n203_ = new_nr_ & new_ns_ & new_na0_;
  assign new_nz1_ = new_nc0_ | new_nd0_;
  assign new_n_n174_ = new_n_n14_ & new_n_n15_ & new_n_n12_ & new_n_n13_ & new_nd_ & new_no_ & new_n_n17_ & new_n_n29_ & new_n_n30_ & new_n_n16_;
  assign new_n_n165_ = new_n_n13_ & new_n_n14_ & new_nd_ & new_n_n12_ & new_nb_ & new_nz0_ & new_nl_ & new_no_ & new_n_n30_ & new_n_n17_ & new_n_n16_ & new_n_n15_;
  assign new_n_n133_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n23_ & new_n_n26_ & new_n_n35_ & new_n_n21_ & new_n_n34_ & new_n_n33_;
  assign new_n_n124_ = new_n_n23_ & new_n_n25_ & new_na_ & new_n_n30_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n115_ = new_n_n31_ & new_n_n32_ & new_nn_ & new_n_n23_ & new_n_n26_ & new_n_n35_ & new_n_n38_ & new_n_n34_ & new_n_n33_;
  assign new_n_n106_ = new_n_n32_ & new_n_n33_ & new_n_n22_ & new_n_n31_ & new_n_n25_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n309_ = new_ne0_ & new_no_ & new_n_n37_ & new_n_n41_ & new_n_n40_ & new_np_;
  assign new_n_n299_ = new_n_n26_ & new_np0_ & new_nv_ & new_n_n37_ & new_n_n41_ & new_n_n6_ & new_n_n19_;
  assign new_n_n278_ = new_np0_ & new_n_n41_ & new_nh_ & new_n_n5_ & new_n_n4_ & new_n_n3_;
  assign new_n_n268_ = new_na_ & new_ne0_;
  assign new_n_n217_ = new_nq0_ & new_n_n41_ & new_n_n24_ & new_ni_ & new_ng_ & new_n_n6_;
  assign new_nv1_ = new_n_n204_ | new_n_n206_ | new_n_n205_ | new_n_n207_;
  assign new_n_n199_ = new_nr0_ & new_n_n38_;
  assign new_nd2_ = new_n_n191_ | new_n_n190_ | new_n_n188_ | new_n_n187_ | new_n_n189_ | new_n_n186_ | new_nz_ | new_ni0_ | new_nh0_ | new_ny_ | new_n_n192_;
  assign new_n_n183_ = new_n_n24_ & new_n_n35_ & new_n_n31_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n132_ = new_n_n22_ & new_n_n31_ & new_n_n28_ & new_n_n23_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n121_ = new_n_n31_ & new_n_n32_ & new_nm_ & new_n_n23_ & new_n_n26_ & new_n_n35_ & new_n_n38_ & new_n_n34_ & new_n_n33_;
  assign new_n_n110_ = new_n_n30_ & new_n_n23_ & new_nn_ & new_n_n28_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n99_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n21_ & new_n_n35_;
  assign new_n_n9_ = ~new_nq0_;
  assign new_ng1_ = new_n_n302_ | new_n_n300_ | new_n_n303_ | new_n_n299_ | new_n_n301_ | new_n_n288_ | new_n_n297_ | new_n_n298_ | new_n_n293_ | new_n_n287_ | new_n_n294_ | new_n_n284_ | new_n_n295_ | new_n_n283_ | new_n_n305_ | new_n_n304_ | new_n_n307_ | new_n_n306_ | new_n_n292_ | new_n_n282_ | new_n_n308_ | new_n_n281_ | new_n_n286_ | new_n_n285_ | new_n_n296_ | new_n_n280_ | new_n_n289_ | new_n_n291_ | new_n_n290_;
  assign new_n_n300_ = new_n_n26_ & new_np0_ & new_n_n7_ & new_ng_ & new_n_n41_ & new_n_n37_ & new_n_n19_;
  assign new_n_n277_ = new_nd0_ & new_n_n36_ & new_n_n41_ & new_nh_ & new_n_n5_ & new_n_n4_ & new_n_n3_;
  assign new_n_n269_ = new_ns0_ & new_nm_;
  assign new_n_n216_ = new_n_n7_ & new_n_n41_ & new_n_n24_ & new_ni_ & new_np0_ & new_ng_;
  assign new_n_n208_ = new_n_n24_ & new_n_n1_ & new_nl_ & new_n_n0_ & new_na0_ & new_n_n41_ & new_n_n38_ & new_nb_ & new_n_n40_ & new_nr_;
  assign new_n_n193_ = new_n_n4_ & new_np_ & new_n_n3_ & new_n_n24_ & new_np0_ & new_n_n41_ & new_n_n8_ & new_n_n5_ & new_n_n40_ & new_no_;
  assign new_n_n192_ = new_n_n41_ & new_nv_ & new_np0_ & new_ni_;
  assign new_n_n184_ = new_n_n35_ & new_n_n31_ & new_n_n34_ & new_n_n30_ & new_n_n26_;
  assign new_n_n131_ = new_n_n23_ & new_n_n31_ & new_n_n28_ & new_n_n30_ & new_n_n21_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n122_ = new_n_n30_ & new_n_n23_ & new_na_ & new_n_n28_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n109_ = new_n_n34_ & new_n_n35_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n38_ & new_n_n21_;
  assign new_n_n100_ = new_n_n25_ & new_n_n31_ & new_n_n30_ & new_n_n23_ & new_n_n29_ & new_nj_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n290_ = new_n_n37_ & new_n_n8_ & new_np0_ & new_n_n19_ & new_n_n40_ & new_n_n24_ & new_n_n7_ & new_n_n41_ & new_n_n25_;
  assign new_nh1_ = new_n_n276_ | new_n_n278_ | new_n_n277_ | new_n_n279_;
  assign new_n_n270_ = new_nq0_ & new_nm_;
  assign new_n_n215_ = new_n_n7_ & new_n_n41_ & new_n_n24_ & new_ni_ & new_ng_ & new_nq0_;
  assign new_n_n201_ = new_ng0_ & new_n_n38_;
  assign new_n_n194_ = new_n_n4_ & new_np_ & new_n_n3_ & new_n_n24_ & new_ne0_ & new_n_n41_ & new_n_n8_ & new_n_n5_ & new_n_n40_ & new_no_;
  assign new_n_n130_ = new_n_n23_ & new_n_n22_ & new_n_n28_ & new_n_n30_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n119_ = new_n_n23_ & new_n_n31_ & new_nm_ & new_n_n30_ & new_n_n38_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n112_ = new_n_n23_ & new_n_n25_ & new_nn_ & new_n_n30_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n101_ = new_n_n31_ & new_n_n32_ & new_n_n23_ & new_n_n25_ & new_n_n29_ & new_n_n26_ & new_n_n35_ & new_nj_ & new_n_n34_ & new_n_n33_;
  assign new_n_n289_ = new_n_n6_ & new_n_n37_ & new_np0_ & new_n_n19_ & new_n_n40_ & new_n_n41_ & new_n_n24_ & new_n_n25_ & new_n_n8_;
  assign new_n_n280_ = new_np0_ & new_n_n6_ & new_n_n1_ & new_n_n36_ & new_n_n40_ & new_n_n41_ & new_n_n24_ & new_n_n8_ & new_n_n37_;
  assign new_n_n279_ = new_ns0_ & new_n_n41_ & new_nh_ & new_n_n5_ & new_n_n4_ & new_n_n3_;
  assign new_n_n207_ = new_n_n41_ & new_n_n40_ & new_n_n38_ & new_n_n24_ & new_ng0_;
  assign new_n_n200_ = new_nf0_ & new_n_n38_;
  assign new_n_n195_ = new_n_n24_ & new_n_n4_ & new_np0_ & new_n_n3_ & new_n_n41_ & new_n_n40_ & new_n_n5_ & new_no_ & new_n_n7_;
  assign new_n_n129_ = new_n_n31_ & new_n_n32_ & new_n_n24_ & new_n_n23_ & new_n_n26_ & new_n_n35_ & new_n_n38_ & new_n_n34_ & new_n_n33_;
  assign new_n_n120_ = new_n_n25_ & new_n_n31_ & new_nm_ & new_n_n23_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n111_ = new_n_n23_ & new_n_n31_ & new_nn_ & new_n_n28_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n102_ = new_n_n31_ & new_n_n32_ & new_n_n25_ & new_n_n22_ & new_n_n30_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n333_ = new_n_n22_ & new_na0_;
  assign new_n_n275_ = new_ne0_ & new_nm_;
  assign new_n_n264_ = new_na_ & new_nk0_;
  assign new_n_n253_ = new_na_ & new_nt_ & new_ni0_;
  assign new_n_n243_ = new_nh_ & new_ne_ & new_ne0_;
  assign new_n_n232_ = new_n_n7_ & new_no_ & new_n_n24_ & new_n_n37_ & new_ne_ & new_nd0_ & new_n_n41_ & new_nd_;
  assign new_n_n189_ = new_n_n41_ & new_ni_ & new_ng_ & new_n_n18_ & new_np0_;
  assign new_n_n179_ = new_np_ & new_no_ & new_nq_ & new_n_n35_ & new_n_n31_ & new_n_n34_ & new_n_n30_ & new_n_n24_;
  assign new_n_n169_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n29_ & new_n_n17_ & new_n_n23_ & new_n_n16_ & new_n_n15_;
  assign new_n_n158_ = new_n_n14_ & new_n_n15_ & new_n_n12_ & new_n_n13_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_no_ & new_n_n17_ & new_n_n23_ & new_n_n30_ & new_n_n16_;
  assign new_n_n148_ = new_ns0_ & new_nh_;
  assign new_n_n139_ = new_n_n31_ & new_n_n32_ & new_n_n23_ & new_n_n25_ & new_n_n26_ & new_n_n35_ & new_n_n21_ & new_n_n34_ & new_n_n33_;
  assign new_n_n5_ = ~new_ne_;
  assign new_n_n334_ = new_n_n21_ & new_na0_;
  assign new_n_n274_ = new_ng0_ & new_nm_;
  assign new_n_n265_ = new_na_ & new_np0_;
  assign new_n_n252_ = new_ng0_ & new_na_ & new_n_n38_;
  assign new_n_n244_ = new_nh_ & new_nu_ & new_ne0_;
  assign new_n_n224_ = new_ns0_ & new_n_n3_ & new_n_n41_ & new_n_n40_ & new_n_n37_ & new_n_n5_ & new_n_n4_;
  assign new_n_n188_ = new_nq0_ & new_n_n41_ & new_ni_ & new_ng_ & new_n_n6_ & new_n_n24_;
  assign new_n_n180_ = new_n_n9_ & new_n_n35_ & new_n_n31_ & new_n_n34_ & new_n_n30_ & new_n_n15_;
  assign new_n_n168_ = new_n_n12_ & new_n_n13_ & new_n_n11_ & new_nd_ & new_n_n10_ & new_n_n29_ & new_n_n16_ & new_n_n17_ & new_n_n15_ & new_n_n14_;
  assign new_n_n159_ = new_nd_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_nb_ & new_nz0_ & new_nl_ & new_n_n17_ & new_n_n15_ & new_n_n16_ & new_n_n14_ & new_n_n13_;
  assign new_n_n147_ = new_nb_ & new_n_n21_ & new_na0_;
  assign new_n_n140_ = new_n_n31_ & new_n_n32_ & new_n_n23_ & new_n_n22_ & new_n_n26_ & new_n_n35_ & new_n_n38_ & new_n_n34_ & new_n_n33_;
  assign new_n_n6_ = ~new_nq_;
  assign new_n_n325_ = new_n_n0_ & new_nv_ & new_na0_ & new_nl_ & new_n_n41_ & new_n_n38_ & new_nb_ & new_n_n40_ & new_n_n39_;
  assign new_n_n317_ = new_n_n40_ & new_n_n41_ & new_n_n18_ & new_n_n37_ & new_ne0_;
  assign new_n_n276_ = new_ne0_ & new_n_n18_ & new_n_n41_ & new_nh_ & new_n_n5_ & new_n_n4_ & new_n_n3_;
  assign new_n_n266_ = new_na_ & new_nd0_;
  assign new_n_n251_ = new_nd_ & new_nw_ & new_nd0_ & new_n_n24_;
  assign new_n_n234_ = new_ne0_ & new_n_n24_ & new_n_n37_ & new_n_n41_ & new_ne_ & new_no_ & new_n_n7_;
  assign new_n_n225_ = new_nh0_ & new_n_n3_ & new_n_n41_ & new_n_n40_ & new_n_n38_ & new_n_n5_ & new_n_n4_;
  assign new_n_n191_ = new_n_n41_ & new_ni_ & new_ng_ & new_n_n6_ & new_np0_;
  assign new_n_n181_ = new_n_n15_ & new_n_n35_ & new_n_n31_ & new_n_n34_ & new_n_n30_ & new_nv_;
  assign new_n_n167_ = new_n_n38_ & new_nb_ & new_n_n40_ & new_nl_ & new_nr_ & new_n_n17_ & new_n_n14_ & new_n_n16_ & new_n_n12_ & new_n_n37_;
  assign new_n_n156_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_n_n23_ & new_n_n30_ & new_n_n17_ & new_n_n16_ & new_n_n15_;
  assign new_n_n150_ = new_na0_ & new_n_n22_;
  assign new_n_n141_ = new_n_n32_ & new_n_n33_ & new_n_n23_ & new_n_n31_ & new_n_n26_ & new_n_n21_ & new_n_n38_ & new_n_n35_ & new_n_n34_;
  assign new_n_n7_ = ~new_np_;
  assign new_nc1_ = new_n_n323_ | new_n_n324_;
  assign new_n_n318_ = new_nu0_ & new_no0_;
  assign new_nk1_ = new_n_n268_ | new_n_n264_ | new_n_n266_ | new_n_n269_ | new_n_n267_ | new_n_n270_ | new_n_n255_ | new_n_n254_ | new_n_n265_ | new_n_n260_ | new_n_n261_ | new_n_n251_ | new_n_n262_ | new_n_n263_ | new_n_n253_ | new_n_n252_ | new_n_n257_ | new_n_n256_ | new_n_n272_ | new_n_n271_ | new_n_n274_ | new_n_n273_ | new_n_n258_ | new_n_n275_ | new_n_n259_;
  assign new_n_n267_ = new_na_ & new_nh0_;
  assign new_n_n242_ = new_nb_ & new_nk_ & new_na0_;
  assign new_n_n233_ = new_n_n7_ & new_no_ & new_n_n24_ & new_n_n37_ & new_nd0_ & new_nu_ & new_n_n41_ & new_nd_;
  assign new_n_n226_ = new_n_n40_ & new_n_n41_ & new_ng0_ & new_nj_ & new_n_n25_ & new_n_n37_;
  assign new_n_n190_ = new_n_n41_ & new_ni_ & new_ng_ & new_n_n7_ & new_np0_;
  assign new_n_n182_ = new_n_n15_ & new_n_n35_ & new_n_n31_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n166_ = new_n_n14_ & new_n_n15_ & new_n_n12_ & new_n_n13_ & new_nb_ & new_nz0_ & new_nl_ & new_no_ & new_n_n17_ & new_n_n23_ & new_n_n30_ & new_n_n16_;
  assign new_n_n157_ = new_n_n13_ & new_n_n14_ & new_nd_ & new_n_n12_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_no_ & new_n_n30_ & new_n_n17_ & new_n_n16_ & new_n_n15_;
  assign new_n_n149_ = new_np0_ & new_nh_;
  assign new_nh2_ = new_n_n136_ | new_n_n135_ | new_n_n133_ | new_n_n132_ | new_n_n134_ | new_n_n82_ | new_n_n64_ | new_n_n73_ | new_n_n55_ | new_n_n72_ | new_n_n83_ | new_n_n65_ | new_n_n84_ | new_n_n54_ | new_n_n75_ | new_n_n53_ | new_n_n62_ | new_n_n85_ | new_n_n63_ | new_n_n74_ | new_n_n52_ | new_n_n121_ | new_n_n130_ | new_n_n77_ | new_n_n86_ | new_n_n68_ | new_n_n131_ | new_n_n59_ | new_n_n120_ | new_n_n76_ | new_n_n87_ | new_n_n69_ | new_n_n110_ | new_n_n58_ | new_n_n101_ | new_n_n79_ | new_n_n88_ | new_n_n66_ | new_n_n111_ | new_n_n57_ | new_n_n100_ | new_n_n78_ | new_n_n89_ | new_n_n67_ | new_n_n126_ | new_n_n56_ | new_n_n108_ | new_n_n117_ | new_n_n99_ | new_n_n81_ | new_n_n90_ | new_n_n127_ | new_n_n109_ | new_n_n116_ | new_n_n98_ | new_n_n80_ | new_n_n91_ | new_n_n128_ | new_n_n106_ | new_n_n119_ | new_n_n97_ | new_n_n61_ | new_n_n70_ | new_n_n129_ | new_n_n107_ | new_n_n118_ | new_n_n96_ | new_n_n60_ | new_n_n71_ | new_n_n113_ | new_n_n122_ | new_n_n104_ | new_n_n50_ | new_n_n95_ | new_n_n94_ | new_n_n124_ | new_n_n51_ | new_n_n123_ | new_n_n105_ | new_n_n112_ | new_n_n92_ | new_n_n139_ | new_n_n141_ | new_n_n140_ | new_n_n138_ | new_n_n137_ | new_n_n125_ | new_n_n103_ | new_n_n114_ | new_n_n115_ | new_n_n93_ | new_n_n102_;
  assign new_n_n8_ = ~new_ng_;
  assign new_na1_ = new_n_n333_ | new_n_n332_ | new_n_n335_ | new_n_n334_ | new_n_n330_ | new_n_n336_ | new_n_n331_;
  assign new_n_n327_ = new_nk0_ & new_nv_ & new_n_n41_ & new_n_n38_ & new_nb_ & new_n_n40_ & new_n_n39_;
  assign new_ne1_ = new_n_n316_ | new_n_n318_ | new_n_n317_ | new_n_n315_ | new_n_n314_;
  assign new_n_n316_ = new_nd0_ & new_nd_ & new_n_n40_ & new_ng_ & new_n_n18_ & new_nu_;
  assign new_n_n307_ = new_nv0_ & new_no0_;
  assign new_n_n296_ = new_n_n1_ & new_n_n26_ & new_n_n7_ & new_n_n41_ & new_nv_ & new_n_n37_ & new_np0_;
  assign new_n_n285_ = new_n_n37_ & new_n_n8_ & new_n_n1_ & new_np0_ & new_n_n40_ & new_n_n24_ & new_n_n18_ & new_n_n41_ & new_n_n25_;
  assign new_n_n271_ = new_nk0_ & new_nm_;
  assign new_n_n257_ = new_nm_ & new_n_n24_ & new_nc0_;
  assign new_n_n247_ = new_nf0_ & new_nb_;
  assign new_n_n236_ = new_n_n24_ & new_n_n8_ & new_n_n37_ & new_ne_ & new_nd0_ & new_n_n41_ & new_nd_;
  assign new_n_n227_ = new_n_n41_ & new_n_n38_ & new_nf_ & new_nv_ & new_ng0_;
  assign new_n_n214_ = new_n_n18_ & new_n_n41_ & new_n_n24_ & new_ni_ & new_np0_ & new_ng_;
  assign new_n_n205_ = new_n_n19_ & new_n_n41_ & new_n_n40_ & new_n_n38_ & new_n_n24_ & new_nk0_;
  assign new_n_n197_ = new_n_n34_ & new_n_n17_ & new_n_n31_ & new_n_n28_ & new_n_n14_;
  assign new_ne2_ = new_n_n182_ | new_n_n181_ | new_n_n184_ | new_n_n183_ | new_n_n180_ | new_n_n179_ | new_n_n185_ | new_n_n178_;
  assign new_n_n176_ = new_nl_ & new_nb_ & new_nz0_ & new_n_n17_ & new_n_n14_ & new_n_n16_ & new_n_n12_ & new_n_n37_;
  assign new_n_n173_ = new_n_n14_ & new_n_n15_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n29_ & new_n_n17_ & new_n_n23_ & new_n_n30_ & new_n_n16_;
  assign new_n_n162_ = new_n_n13_ & new_n_n14_ & new_n_n10_ & new_n_n12_ & new_nb_ & new_nz0_ & new_nl_ & new_no_ & new_n_n17_ & new_n_n23_ & new_n_n16_ & new_n_n15_;
  assign new_n_n151_ = new_nd_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_n_n17_ & new_n_n15_ & new_n_n16_ & new_n_n14_ & new_n_n13_;
  assign new_n_n142_ = new_nb_ & new_n_n20_ & new_nj_ & new_na0_;
  assign new_n_n118_ = new_n_n23_ & new_n_n25_ & new_nm_ & new_n_n30_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n107_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n25_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n21_ & new_n_n35_;
  assign new_n_n1_ = ~new_ns_;
  assign new_n_n326_ = new_nl_ & new_n_n0_ & new_na0_ & new_n_n41_ & new_nj_ & new_nb_ & new_n_n40_ & new_n_n39_;
  assign new_n_n319_ = new_n_n18_ & new_nd0_ & new_n_n24_ & new_n_n41_ & new_n_n40_ & new_n_n36_ & new_n_n37_;
  assign new_n_n315_ = new_ne_ & new_nd_ & new_n_n40_ & new_ng_ & new_n_n18_ & new_nd0_;
  assign new_n_n308_ = new_nd0_ & new_nv_;
  assign new_n_n295_ = new_n_n1_ & new_n_n26_ & new_n_n18_ & new_ng_ & new_n_n41_ & new_n_n37_ & new_np0_;
  assign new_n_n286_ = new_n_n19_ & new_n_n6_ & new_n_n36_ & new_np0_ & new_n_n40_ & new_n_n41_ & new_n_n24_ & new_n_n8_ & new_n_n37_;
  assign new_n_n261_ = new_na0_ & new_na_;
  assign new_n_n256_ = new_nm_ & new_n_n24_ & new_nb0_;
  assign new_n_n248_ = new_nw_ & new_nh0_;
  assign new_n_n235_ = new_ne0_ & new_n_n24_ & new_n_n37_ & new_n_n41_ & new_nu_ & new_no_ & new_n_n7_;
  assign new_nn1_ = new_n_n224_ | new_n_n223_ | new_n_n226_ | new_n_n225_ | new_n_n222_ | new_n_n221_ | new_n_n227_ | new_n_n220_;
  assign new_n_n223_ = new_nw0_ & new_no0_ & new_n_n41_ & new_n_n5_ & new_n_n40_ & new_n_n4_ & new_n_n3_;
  assign new_n_n204_ = new_n_n2_ & new_n_n41_ & new_n_n40_ & new_n_n38_ & new_nv_ & new_ng0_;
  assign new_n_n198_ = new_nj_ & new_n_n34_ & new_n_n31_;
  assign new_n_n185_ = new_na_ & new_n_n34_ & new_n_n35_ & new_n_n31_ & new_n_n30_;
  assign new_n_n177_ = new_n_n37_ & new_n_n29_ & new_n_n16_ & new_n_n17_ & new_n_n14_ & new_n_n12_;
  assign new_n_n172_ = new_n_n13_ & new_n_n14_ & new_nd_ & new_n_n12_ & new_n_n11_ & new_n_n29_ & new_n_n30_ & new_n_n17_ & new_n_n16_ & new_n_n15_;
  assign new_n_n163_ = new_n_n12_ & new_n_n13_ & new_n_n11_ & new_nd_ & new_nb_ & new_nz0_ & new_nl_ & new_n_n17_ & new_n_n16_ & new_n_n30_ & new_n_n15_ & new_n_n14_;
  assign new_ng2_ = new_nm0_ | new_n_n150_ | new_nr0_ | new_nx0_ | new_n_n142_ | new_nf0_ | new_n_n143_ | new_n_n148_ | new_ns1_ | new_n_n149_ | new_n_n146_ | new_n_n147_ | new_n_n145_ | new_n_n144_;
  assign new_n_n143_ = new_nb_ & new_n_n20_ & new_nm_ & new_na0_;
  assign new_n_n117_ = new_n_n23_ & new_n_n31_ & new_nm_ & new_n_n28_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n108_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n22_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n38_ & new_n_n35_;
  assign new_n_n2_ = ~new_nf_;
  assign new_n_n335_ = new_nm_ & new_na0_;
  assign new_n_n329_ = new_nt0_ & new_no0_;
  assign new_n_n320_ = new_nd0_ & new_n_n7_ & new_n_n24_ & new_n_n41_ & new_n_n40_ & new_n_n36_ & new_n_n37_;
  assign new_n_n314_ = new_n_n3_ & new_n_n5_ & new_nd_ & new_n_n18_ & new_n_n40_ & new_n_n4_ & new_nd0_;
  assign new_n_n305_ = new_ng_ & new_nd0_ & new_ne_ & new_no_ & new_n_n40_ & new_np_ & new_n_n24_;
  assign new_n_n298_ = new_n_n26_ & new_np0_ & new_n_n41_ & new_n_n37_ & new_ng_ & new_n_n6_ & new_n_n19_;
  assign new_n_n287_ = new_n_n19_ & new_n_n37_ & new_n_n36_ & new_np0_ & new_n_n40_ & new_n_n24_ & new_n_n7_ & new_n_n41_ & new_n_n8_;
  assign new_n_n273_ = new_nh0_ & new_nm_;
  assign new_n_n262_ = new_na_ & new_ns0_;
  assign new_n_n255_ = new_np0_ & new_nr_ & new_ns_;
  assign new_n_n245_ = new_nh_ & new_nd0_ & new_ne_;
  assign new_n_n238_ = new_ne0_ & new_n_n37_ & new_n_n41_ & new_ne_ & new_n_n8_ & new_n_n24_;
  assign new_n_n228_ = new_n_n4_ & new_n_n7_ & new_n_n3_ & new_n_n24_ & new_nd0_ & new_n_n41_ & new_n_n5_ & new_nd_ & new_n_n40_ & new_no_;
  assign new_n_n222_ = new_n_n3_ & new_n_n4_ & new_ne0_ & new_n_n41_ & new_n_n5_ & new_n_n40_ & new_no_ & new_n_n7_;
  assign new_nr1_ = new_n_n210_ | new_n_n212_ | new_n_n211_ | new_n_n209_ | new_n_n208_;
  assign new_ny1_ = new_n_n197_ | new_n_n198_;
  assign new_n_n187_ = new_n_n7_ & new_n_n41_ & new_ni_ & new_ng_ & new_n_n24_ & new_nq0_;
  assign new_nf2_ = new_n_n174_ | new_n_n173_ | new_n_n176_ | new_n_n175_ | new_n_n151_ | new_n_n177_ | new_n_n161_ | new_n_n164_ | new_n_n165_ | new_n_n155_ | new_n_n158_ | new_n_n154_ | new_n_n160_ | new_n_n159_ | new_n_n171_ | new_n_n169_ | new_n_n172_ | new_n_n170_ | new_n_n166_ | new_n_n168_ | new_n_n157_ | new_n_n156_ | new_n_n167_ | new_n_n153_ | new_n_n162_ | new_n_n152_ | new_n_n163_;
  assign new_n_n171_ = new_n_n14_ & new_n_n15_ & new_n_n12_ & new_n_n13_ & new_n_n10_ & new_no_ & new_n_n23_ & new_n_n29_ & new_n_n17_ & new_n_n16_;
  assign new_n_n160_ = new_n_n12_ & new_n_n13_ & new_n_n10_ & new_n_n11_ & new_nb_ & new_nz0_ & new_nl_ & new_n_n23_ & new_n_n16_ & new_n_n17_ & new_n_n15_ & new_n_n14_;
  assign new_n_n153_ = new_n_n12_ & new_n_n13_ & new_n_n10_ & new_nd_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_no_ & new_n_n16_ & new_n_n17_ & new_n_n15_ & new_n_n14_;
  assign new_n_n144_ = new_nb_ & new_n_n19_ & new_n_n20_ & new_na0_;
  assign new_n_n138_ = new_n_n22_ & new_n_n31_ & new_n_n23_ & new_n_n25_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n127_ = new_n_n31_ & new_n_n32_ & new_na_ & new_n_n23_ & new_n_n26_ & new_n_n35_ & new_n_n38_ & new_n_n34_ & new_n_n33_;
  assign new_n_n3_ = ~new_nw_;
  assign new_n_n336_ = new_nn_ & new_na0_;
  assign new_n_n328_ = new_nj_ & new_n_n3_ & new_ng0_ & new_nc_;
  assign new_n_n321_ = new_n_n24_ & new_nc0_ & new_n_n40_;
  assign new_nf1_ = new_n_n311_ | new_n_n313_ | new_n_n312_ | new_n_n310_ | new_n_n309_;
  assign new_n_n306_ = new_nd0_ & new_n_n24_ & new_n_n5_ & new_no_ & new_n_n40_ & new_np_ & new_n_n4_;
  assign new_n_n297_ = new_n_n1_ & new_n_n26_ & new_n_n18_ & new_n_n41_ & new_nv_ & new_n_n37_ & new_np0_;
  assign new_n_n288_ = new_n_n19_ & new_n_n37_ & new_n_n36_ & new_np0_ & new_n_n40_ & new_n_n24_ & new_n_n18_ & new_n_n41_ & new_n_n8_;
  assign new_n_n272_ = new_nr0_ & new_nb_;
  assign new_n_n263_ = new_na_ & new_nq0_;
  assign new_n_n254_ = new_nr_ & new_ns_ & new_nl0_;
  assign new_n_n246_ = new_nh_ & new_nu_ & new_nd0_;
  assign new_n_n237_ = new_n_n24_ & new_n_n8_ & new_n_n37_ & new_nd0_ & new_nu_ & new_n_n41_ & new_nd_;
  assign new_n_n229_ = new_nh0_ & new_nj_;
  assign new_n_n221_ = new_n_n3_ & new_n_n4_ & new_n_n6_ & new_n_n8_ & new_nq0_ & new_n_n41_ & new_n_n5_ & new_n_n40_ & new_no_ & new_np_;
  assign new_n_n213_ = new_n_n18_ & new_n_n41_ & new_n_n24_ & new_ni_ & new_ng_ & new_nq0_;
  assign new_n_n206_ = new_nk0_ & new_n_n41_ & new_n_n40_ & new_n_n38_ & new_nn_ & new_nv_;
  assign new_n_n186_ = new_n_n18_ & new_n_n41_ & new_ni_ & new_ng_ & new_n_n24_ & new_nq0_;
  assign new_n_n178_ = new_np_ & new_no_ & new_nq_ & new_n_n35_ & new_n_n31_ & new_n_n34_ & new_n_n30_ & new_n_n15_;
  assign new_n_n170_ = new_n_n13_ & new_n_n14_ & new_nd_ & new_n_n12_ & new_n_n10_ & new_no_ & new_n_n17_ & new_n_n29_ & new_n_n16_ & new_n_n15_;
  assign new_n_n161_ = new_n_n12_ & new_n_n13_ & new_n_n10_ & new_nd_ & new_nb_ & new_nz0_ & new_nl_ & new_no_ & new_n_n16_ & new_n_n17_ & new_n_n15_ & new_n_n14_;
  assign new_n_n152_ = new_n_n12_ & new_n_n13_ & new_n_n10_ & new_n_n11_ & new_nb_ & new_nl_ & new_n_n38_ & new_nr_ & new_n_n40_ & new_n_n23_ & new_n_n16_ & new_n_n17_ & new_n_n15_ & new_n_n14_;
  assign new_n_n145_ = new_nh_ & new_n_n36_ & new_nd0_;
  assign new_n_n137_ = new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n23_ & new_n_n38_ & new_n_n35_ & new_n_n21_ & new_n_n34_ & new_n_n33_;
  assign new_n_n128_ = new_n_n23_ & new_n_n31_ & new_n_n24_ & new_n_n30_ & new_n_n38_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n4_ = ~new_nu_;
  assign new_n_n93_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n24_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n38_ & new_n_n35_;
  assign new_n_n82_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_na_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n71_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_nn_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n60_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n28_ & new_n_n36_ & new_nj_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_ni2_ = new_n_n48_ | new_n_n46_ | new_n_n49_ | new_n_n47_ | new_n_n43_ | new_n_n45_ | new_nb0_ | new_ny_ | new_nh0_ | new_nc0_ | new_n_n44_ | new_nz_ | new_n_n42_;
  assign new_n_n94_ = new_n_n23_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nj_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n81_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_nm_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n38_ & new_n_n35_;
  assign new_n_n72_ = new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n25_ & new_nn_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n59_ = new_n_n32_ & new_n_n33_ & new_n_n25_ & new_n_n31_ & new_n_n29_ & new_n_n24_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n50_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n27_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n95_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n23_ & new_n_n28_ & new_n_n26_ & new_n_n35_ & new_nj_ & new_n_n34_ & new_n_n33_;
  assign new_n_n80_ = new_n_n32_ & new_n_n33_ & new_n_n25_ & new_n_n31_ & new_nm_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n69_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n23_ & new_n_n27_ & new_n_n26_ & new_n_n35_ & new_n_n38_ & new_n_n34_ & new_n_n33_;
  assign new_n_n62_ = new_n_n32_ & new_n_n33_ & new_n_n25_ & new_n_n31_ & new_n_n30_ & new_n_n29_ & new_n_n36_ & new_nj_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n51_ = new_n_n32_ & new_n_n33_ & new_n_n29_ & new_n_n31_ & new_n_n28_ & new_n_n27_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n96_ = new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n22_ & new_n_n28_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n79_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_nm_ & new_n_n36_ & new_n_n38_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n70_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_nn_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n61_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n28_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_nj_ & new_n_n35_;
  assign new_n_n52_ = new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n25_ & new_n_n29_ & new_n_n27_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n0_ = ~new_nk_;
  assign new_n_n97_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n36_ & new_n_n21_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n43_ = new_nv_ & new_n_n39_ & new_nk0_ & new_n_n38_ & new_nb_ & new_n_n41_ & new_nl_ & new_n_n40_;
  assign new_n_n32_ = ~new_nc0_;
  assign new_n_n21_ = ~new_nl_;
  assign new_n_n10_ = ~new_nt_;
  assign new_n_n98_ = new_n_n32_ & new_n_n33_ & new_n_n22_ & new_n_n31_ & new_n_n28_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n42_ = new_n_n39_ & new_n_n40_ & new_nk0_ & new_nv_ & new_nc_ & new_n_n41_ & new_ng0_ & new_nb_ & new_nl_;
  assign new_n_n33_ = ~new_nb0_;
  assign new_n_n20_ = ~new_nz0_;
  assign new_n_n11_ = ~new_ne0_;
  assign new_n_n41_ = ~new_na_;
  assign new_n_n30_ = ~new_ni0_;
  assign new_n_n23_ = ~new_nd0_;
  assign new_n_n12_ = ~new_nx0_;
  assign new_n_n40_ = ~new_nm_;
  assign new_n_n31_ = ~new_nh0_;
  assign new_n_n22_ = ~new_nb_;
  assign new_n_n13_ = ~new_ns0_;
  assign new_n_n68_ = new_n_n25_ & new_n_n31_ & new_n_n29_ & new_n_n23_ & new_n_n27_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n57_ = new_n_n32_ & new_n_n33_ & new_n_n29_ & new_n_n31_ & new_n_n28_ & new_n_n24_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n47_ = new_nd_ & new_nd0_;
  assign new_n_n36_ = ~new_nd_;
  assign new_n_n25_ = ~new_nc_;
  assign new_n_n14_ = ~new_nr0_;
  assign new_n_n67_ = new_n_n23_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n38_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n58_ = new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n25_ & new_n_n29_ & new_n_n24_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n46_ = new_nc_ & new_nj_ & new_ng0_;
  assign new_n_n37_ = ~new_nh_;
  assign new_n_n24_ = ~new_nv_;
  assign new_n_n15_ = ~new_np0_;
  assign new_n_n88_ = new_n_n30_ & new_n_n23_ & new_n_n28_ & new_n_n29_ & new_n_n24_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n77_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_nm_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n45_ = new_na0_ & new_n_n39_ & new_nj_ & new_nb_ & new_n_n41_ & new_nl_ & new_n_n40_;
  assign new_n_n34_ = ~new_nz_;
  assign new_n_n27_ = ~new_nk0_;
  assign new_n_n16_ = ~new_nm0_;
  assign new_n_n87_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_na_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n38_ & new_n_n35_;
  assign new_n_n78_ = new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n25_ & new_nm_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n44_ = new_na0_ & new_nv_ & new_n_n41_ & new_nl_ & new_nb_ & new_n_n40_ & new_n_n39_;
  assign new_n_n35_ = ~new_ny_;
  assign new_n_n26_ = ~new_ni_;
  assign new_n_n17_ = ~new_nf0_;
  assign new_n_n89_ = new_n_n23_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n86_ = new_n_n32_ & new_n_n33_ & new_n_n25_ & new_n_n31_ & new_na_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n75_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_nn_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n38_ & new_n_n35_;
  assign new_n_n64_ = new_n_n30_ & new_n_n23_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n53_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n36_ & new_n_n38_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n29_ = ~new_na0_;
  assign new_n_n18_ = ~new_no_;
  assign new_n_n90_ = new_n_n23_ & new_n_n25_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n85_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_na_ & new_n_n36_ & new_n_n38_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n76_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_nm_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n63_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n25_ & new_n_n29_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_nj_ & new_n_n35_;
  assign new_n_n54_ = new_n_n32_ & new_n_n33_ & new_n_n25_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n28_ = ~new_ng0_;
  assign new_n_n19_ = ~new_nr_;
  assign new_n_n91_ = new_n_n25_ & new_n_n31_ & new_n_n29_ & new_n_n23_ & new_n_n24_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n84_ = new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n25_ & new_na_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n73_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_nn_ & new_n_n36_ & new_n_n38_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n66_ = new_n_n23_ & new_n_n25_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n35_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n55_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n27_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n38_ & new_n_n35_;
  assign new_n_n49_ = new_ni0_ & new_ni_;
  assign new_n_n38_ = ~new_nj_;
  assign new_n_n92_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n24_ & new_n_n36_ & new_n_n38_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n83_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_na_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n74_ = new_n_n32_ & new_n_n33_ & new_n_n25_ & new_n_n31_ & new_nn_ & new_n_n36_ & new_n_n26_ & new_nh_ & new_n_n35_ & new_n_n34_;
  assign new_n_n65_ = new_n_n23_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_n_n26_ & new_n_n34_ & new_n_n35_ & new_n_n33_ & new_n_n32_;
  assign new_n_n56_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n24_ & new_n_n36_ & new_n_n35_ & new_nh_ & new_n_n34_ & new_n_n33_;
  assign new_n_n48_ = new_nd0_ & new_n_n37_;
  assign new_n_n39_ = ~new_nn_;
endmodule


