// Benchmark "top" written by ABC on Fri Mar 31 12:12:23 2023

module top ( 
    pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv56_13_, pv56_22_, pv88_7_,
    pv88_29_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_, pv56_15_,
    pv56_24_, pv88_9_, pv88_18_, pv88_27_, pv9_5_, pv56_30_, pv88_2_,
    pv88_15_, pv88_26_, pv9_6_, pv24_10_, pv56_31_, pv88_3_, pv88_16_,
    pv88_25_, pv9_7_, pv9_10_, pv56_10_, pv56_21_, pv88_4_, pv88_13_,
    pv88_24_, pv9_8_, pv56_11_, pv56_20_, pv88_5_, pv88_14_, pv88_23_,
    pv56_5_, pv88_11_, pv88_22_, pv56_4_, pv88_12_, pv88_21_, pv56_7_,
    pv88_20_, pv56_6_, pv88_10_, pv24_8_, pv56_9_, pv24_9_, pv56_8_,
    pv24_6_, pv24_7_, pv24_4_, pv24_5_, pv24_2_, pv24_3_, pv24_0_, pv56_1_,
    pv24_1_, pv56_0_, pv88_30_, pv56_3_, pv88_31_, pv56_2_, pv9_1_,
    pv24_13_, pv9_2_, pv24_14_, pv9_3_, pv24_11_, pv88_0_, pv24_12_,
    pv88_1_, pv56_16_, pv56_27_, pv56_17_, pv56_26_, pv56_18_, pv56_29_,
    pv9_0_, pv56_19_, pv56_28_,
    pv119_1_, pv119_0_, pv119_3_, pv119_30_, pv119_2_, pv151_1_, pv151_18_,
    pv151_0_, pv151_19_, pv119_21_, pv151_3_, pv151_16_, pv119_20_,
    pv151_2_, pv151_17_, pv119_9_, pv119_23_, pv151_27_, pv119_8_,
    pv119_22_, pv151_26_, pv119_25_, pv151_29_, pv119_24_, pv151_28_,
    pv119_5_, pv119_27_, pv119_4_, pv119_26_, pv119_7_, pv119_29_,
    pv119_6_, pv119_28_, pv119_18_, pv119_19_, pv119_16_, pv151_21_,
    pv119_17_, pv151_20_, pv119_14_, pv151_23_, pv119_15_, pv151_22_,
    pv119_12_, pv151_25_, pv151_30_, pv119_13_, pv151_24_, pv151_31_,
    pv119_10_, pv151_5_, pv151_14_, pv119_11_, pv151_4_, pv151_15_,
    pv151_7_, pv151_12_, pv151_6_, pv151_13_, pv151_9_, pv151_10_,
    pv151_8_, pv151_11_  );
  input  pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv56_13_, pv56_22_,
    pv88_7_, pv88_29_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_,
    pv56_15_, pv56_24_, pv88_9_, pv88_18_, pv88_27_, pv9_5_, pv56_30_,
    pv88_2_, pv88_15_, pv88_26_, pv9_6_, pv24_10_, pv56_31_, pv88_3_,
    pv88_16_, pv88_25_, pv9_7_, pv9_10_, pv56_10_, pv56_21_, pv88_4_,
    pv88_13_, pv88_24_, pv9_8_, pv56_11_, pv56_20_, pv88_5_, pv88_14_,
    pv88_23_, pv56_5_, pv88_11_, pv88_22_, pv56_4_, pv88_12_, pv88_21_,
    pv56_7_, pv88_20_, pv56_6_, pv88_10_, pv24_8_, pv56_9_, pv24_9_,
    pv56_8_, pv24_6_, pv24_7_, pv24_4_, pv24_5_, pv24_2_, pv24_3_, pv24_0_,
    pv56_1_, pv24_1_, pv56_0_, pv88_30_, pv56_3_, pv88_31_, pv56_2_,
    pv9_1_, pv24_13_, pv9_2_, pv24_14_, pv9_3_, pv24_11_, pv88_0_,
    pv24_12_, pv88_1_, pv56_16_, pv56_27_, pv56_17_, pv56_26_, pv56_18_,
    pv56_29_, pv9_0_, pv56_19_, pv56_28_;
  output pv119_1_, pv119_0_, pv119_3_, pv119_30_, pv119_2_, pv151_1_,
    pv151_18_, pv151_0_, pv151_19_, pv119_21_, pv151_3_, pv151_16_,
    pv119_20_, pv151_2_, pv151_17_, pv119_9_, pv119_23_, pv151_27_,
    pv119_8_, pv119_22_, pv151_26_, pv119_25_, pv151_29_, pv119_24_,
    pv151_28_, pv119_5_, pv119_27_, pv119_4_, pv119_26_, pv119_7_,
    pv119_29_, pv119_6_, pv119_28_, pv119_18_, pv119_19_, pv119_16_,
    pv151_21_, pv119_17_, pv151_20_, pv119_14_, pv151_23_, pv119_15_,
    pv151_22_, pv119_12_, pv151_25_, pv151_30_, pv119_13_, pv151_24_,
    pv151_31_, pv119_10_, pv151_5_, pv151_14_, pv119_11_, pv151_4_,
    pv151_15_, pv151_7_, pv151_12_, pv151_6_, pv151_13_, pv151_9_,
    pv151_10_, pv151_8_, pv151_11_;
  wire new_n_n127_, new_n_n138_, new_n_n109_, new_n_n76_, new_n_n128_,
    new_n_n137_, new_n_n110_, new_n_n86_, new_n_n129_, new_n_n140_,
    new_n_n111_, new_n_n74_, new_n_n85_, new_n_n130_, new_n_n139_,
    new_n_n112_, new_n_n75_, new_n_n84_, new_n_n150_, new_n_n145_,
    new_n_n105_, new_n_n72_, new_n_n83_, new_n_n149_, new_n_n99_,
    new_n_n146_, new_n_n106_, new_n_n73_, new_n_n82_, new_n_n148_,
    new_n_n152_, new_n_n125_, new_n_n136_, new_n_n107_, new_n_n70_,
    new_n_n81_, new_n_n147_, new_n_n126_, new_n_n135_, new_n_n108_,
    new_n_n71_, new_n_n80_, new_n_n120_, new_n_n114_, new_n_n79_,
    new_n_n119_, new_n_n69_, new_n_n78_, new_n_n122_, new_n_n77_,
    new_n_n121_, new_n_n113_, new_n_n97_, new_n_n124_, new_n_n98_,
    new_n_n123_, new_n_n95_, new_n_n96_, new_n_n93_, new_n_n94_,
    new_n_n91_, new_n_n92_, new_n_n89_, new_n_n116_, new_n_n90_,
    new_n_n115_, new_n_n87_, new_n_n118_, new_n_n88_, new_n_n117_,
    new_n_n154_, new_n_n102_, new_n_n153_, new_n_n103_, new_n_n155_,
    new_n_n100_, new_n_n68_, new_n_n101_, new_n_n104_, new_n_n131_,
    new_n_n142_, new_n_n132_, new_n_n141_, new_n_n133_, new_n_n144_,
    new_n_n151_, new_n_n134_, new_n_n143_, new_nv158_, new_n_n3_,
    new_n_n63_, new_nv197_, new_n_n41_, new_nv210_, new_nv221_, new_nv232_,
    new_nv243_, new_nv265_, new_n_n21_, new_n_n10_, new_nv303_, new_nv314_,
    new_nv325_, new_nv336_, new_nv154_, new_n_n2_, new_nv180_, new_nv192_,
    new_nv203_, new_nv209_, new_nv222_, new_nv231_, new_nv244_, new_nv264_,
    new_n_n20_, new_n_n11_, new_nv304_, new_nv313_, new_nv326_, new_nv335_,
    new_nv162_, new_nv171_, new_n_n64_, new_n_n51_, new_nv198_, new_nv208_,
    new_nv223_, new_nv234_, new_nv241_, new_nv263_, new_nv289_, new_n_n30_,
    new_nv305_, new_nv316_, new_nv323_, new_nv334_, new_nv161_, new_n_n4_,
    new_nv179_, new_nv193_, new_n_n46_, new_nv202_, new_nv224_, new_nv233_,
    new_nv242_, new_nv251_, new_nv290_, new_n_n31_, new_nv306_, new_nv315_,
    new_nv324_, new_nv333_, new_nv165_, new_n_n61_, new_nv188_, new_nv225_,
    new_nv236_, new_nv247_, new_nv269_, new_nv280_, new_nv307_, new_nv318_,
    new_nv329_, new_nv340_, new_nv441_, new_nv163_, new_nv183_, new_n_n56_,
    new_nv226_, new_nv235_, new_nv268_, new_nv270_, new_nv279_, new_nv308_,
    new_nv317_, new_nv330_, new_nv339_, new_nv176_, new_n_n62_, new_nv187_,
    new_nv227_, new_nv245_, new_nv267_, new_nv309_, new_nv320_, new_nv327_,
    new_nv338_, new_n_n67_, new_nv181_, new_nv182_, new_nv237_, new_nv246_,
    new_nv266_, new_nv310_, new_nv319_, new_nv328_, new_nv337_, new_n_n59_,
    new_nv190_, new_n_n48_, new_nv201_, new_n_n37_, new_nv273_, new_nv284_,
    new_n_n35_, new_n_n24_, new_n_n13_, new_nv300_, new_nv164_, new_nv185_,
    new_n_n54_, new_nv196_, new_n_n43_, new_nv217_, new_nv274_, new_nv283_,
    new_n_n34_, new_n_n25_, new_n_n12_, new_nv299_, new_nv166_, new_n_n60_,
    new_nv189_, new_n_n47_, new_n_n38_, new_nv216_, new_nv271_, new_nv282_,
    new_n_n33_, new_n_n22_, new_n_n15_, new_nv298_, new_nv437_, new_nv184_,
    new_n_n55_, new_n_n42_, new_nv206_, new_nv215_, new_nv272_, new_nv281_,
    new_n_n32_, new_n_n23_, new_n_n14_, new_n_n5_, new_nv440_, new_nv169_,
    new_n_n65_, new_n_n57_, new_n_n50_, new_nv199_, new_n_n39_, new_nv214_,
    new_nv228_, new_nv239_, new_nv250_, new_nv277_, new_nv288_, new_nv291_,
    new_n_n28_, new_n_n17_, new_n_n6_, new_nv321_, new_nv332_, new_nv156_,
    new_nv170_, new_nv178_, new_n_n52_, new_nv194_, new_n_n45_, new_nv205_,
    new_nv213_, new_nv218_, new_nv240_, new_nv249_, new_nv278_, new_nv287_,
    new_nv292_, new_n_n29_, new_n_n16_, new_n_n7_, new_nv322_, new_nv331_,
    new_nv157_, new_nv153_, new_nv167_, new_n_n66_, new_n_n58_, new_nv191_,
    new_n_n49_, new_nv200_, new_n_n40_, new_nv212_, new_nv219_, new_nv230_,
    new_nv248_, new_nv275_, new_nv286_, new_nv293_, new_n_n26_, new_n_n19_,
    new_n_n8_, new_nv301_, new_nv312_, new_nv159_, new_nv152_, new_nv168_,
    new_nv177_, new_nv186_, new_n_n53_, new_nv195_, new_n_n44_, new_nv204_,
    new_nv211_, new_nv220_, new_nv229_, new_nv238_, new_nv276_, new_nv285_,
    new_n_n36_, new_n_n27_, new_n_n18_, new_n_n9_, new_nv302_, new_nv311_,
    new_nv160_, new_nv346_, new_nv357_, new_nv368_, new_nv379_, new_nv390_,
    new_nv345_, new_nv358_, new_nv367_, new_nv380_, new_nv389_, new_nv344_,
    new_nv359_, new_nv370_, new_nv377_, new_nv388_, new_nv343_, new_nv360_,
    new_nv369_, new_nv378_, new_nv387_, new_nv155_, new_nv342_, new_nv397_,
    new_nv408_, new_nv419_, new_nv297_, new_nv341_, new_nv398_, new_nv407_,
    new_nv420_, new_nv296_, new_nv399_, new_nv410_, new_nv417_, new_nv295_,
    new_nv400_, new_nv409_, new_nv418_, new_nv294_, new_nv371_, new_nv382_,
    new_nv393_, new_nv404_, new_nv415_, new_nv207_, new_nv372_, new_nv381_,
    new_nv394_, new_nv403_, new_nv416_, new_nv425_, new_nv351_, new_nv362_,
    new_nv395_, new_nv406_, new_nv413_, new_nv424_, new_nv352_, new_nv361_,
    new_nv396_, new_nv405_, new_nv414_, new_nv423_, new_nv350_, new_nv353_,
    new_nv364_, new_nv375_, new_nv386_, new_nv411_, new_nv422_, new_nv349_,
    new_nv354_, new_nv363_, new_nv376_, new_nv385_, new_nv412_, new_nv421_,
    new_nv348_, new_nv355_, new_nv366_, new_nv373_, new_nv384_, new_nv391_,
    new_nv402_, new_nv347_, new_nv356_, new_nv365_, new_nv374_, new_nv383_,
    new_nv392_, new_nv401_;
  assign new_n_n127_ = pv56_12_;
  assign new_n_n138_ = pv56_23_;
  assign new_n_n109_ = pv88_6_;
  assign new_n_n76_ = pv88_19_;
  assign pv119_1_ = new_n_n38_;
  assign new_n_n128_ = pv56_13_;
  assign new_n_n137_ = pv56_22_;
  assign new_n_n110_ = pv88_7_;
  assign new_n_n86_ = pv88_29_;
  assign pv119_0_ = new_n_n37_;
  assign new_n_n129_ = pv56_14_;
  assign new_n_n140_ = pv56_25_;
  assign new_n_n111_ = pv88_8_;
  assign new_n_n74_ = pv88_17_;
  assign new_n_n85_ = pv88_28_;
  assign pv119_3_ = new_n_n40_;
  assign pv119_30_ = new_n_n67_;
  assign new_n_n130_ = pv56_15_;
  assign new_n_n139_ = pv56_24_;
  assign new_n_n112_ = pv88_9_;
  assign new_n_n75_ = pv88_18_;
  assign new_n_n84_ = pv88_27_;
  assign pv119_2_ = new_n_n39_;
  assign new_n_n150_ = pv9_5_;
  assign new_n_n145_ = pv56_30_;
  assign new_n_n105_ = pv88_2_;
  assign new_n_n72_ = pv88_15_;
  assign new_n_n83_ = pv88_26_;
  assign pv151_1_ = new_n_n22_;
  assign pv151_18_ = new_n_n7_;
  assign new_n_n149_ = pv9_6_;
  assign new_n_n99_ = pv24_10_;
  assign new_n_n146_ = pv56_31_;
  assign new_n_n106_ = pv88_3_;
  assign new_n_n73_ = pv88_16_;
  assign new_n_n82_ = pv88_25_;
  assign pv151_0_ = new_n_n21_;
  assign pv151_19_ = new_n_n8_;
  assign new_n_n148_ = pv9_7_;
  assign new_n_n152_ = pv9_10_;
  assign new_n_n125_ = pv56_10_;
  assign new_n_n136_ = pv56_21_;
  assign new_n_n107_ = pv88_4_;
  assign new_n_n70_ = pv88_13_;
  assign new_n_n81_ = pv88_24_;
  assign pv119_21_ = new_n_n58_;
  assign pv151_3_ = new_n_n24_;
  assign pv151_16_ = new_n_n5_;
  assign new_n_n147_ = pv9_8_;
  assign new_n_n126_ = pv56_11_;
  assign new_n_n135_ = pv56_20_;
  assign new_n_n108_ = pv88_5_;
  assign new_n_n71_ = pv88_14_;
  assign new_n_n80_ = pv88_23_;
  assign pv119_20_ = new_n_n57_;
  assign pv151_2_ = new_n_n23_;
  assign pv151_17_ = new_n_n6_;
  assign new_n_n120_ = pv56_5_;
  assign new_n_n114_ = pv88_11_;
  assign new_n_n79_ = pv88_22_;
  assign pv119_9_ = new_n_n46_;
  assign pv119_23_ = new_n_n60_;
  assign pv151_27_ = new_n_n16_;
  assign new_n_n119_ = pv56_4_;
  assign new_n_n69_ = pv88_12_;
  assign new_n_n78_ = pv88_21_;
  assign pv119_8_ = new_n_n45_;
  assign pv119_22_ = new_n_n59_;
  assign pv151_26_ = new_n_n15_;
  assign new_n_n122_ = pv56_7_;
  assign new_n_n77_ = pv88_20_;
  assign pv119_25_ = new_n_n62_;
  assign pv151_29_ = new_n_n18_;
  assign new_n_n121_ = pv56_6_;
  assign new_n_n113_ = pv88_10_;
  assign pv119_24_ = new_n_n61_;
  assign pv151_28_ = new_n_n17_;
  assign new_n_n97_ = pv24_8_;
  assign new_n_n124_ = pv56_9_;
  assign pv119_5_ = new_n_n42_;
  assign pv119_27_ = new_n_n64_;
  assign new_n_n98_ = pv24_9_;
  assign new_n_n123_ = pv56_8_;
  assign pv119_4_ = new_n_n41_;
  assign pv119_26_ = new_n_n63_;
  assign new_n_n95_ = pv24_6_;
  assign pv119_7_ = new_n_n44_;
  assign pv119_29_ = new_n_n66_;
  assign new_n_n96_ = pv24_7_;
  assign pv119_6_ = new_n_n43_;
  assign pv119_28_ = new_n_n65_;
  assign new_n_n93_ = pv24_4_;
  assign pv119_18_ = new_n_n55_;
  assign new_n_n94_ = pv24_5_;
  assign pv119_19_ = new_n_n56_;
  assign new_n_n91_ = pv24_2_;
  assign pv119_16_ = new_n_n53_;
  assign pv151_21_ = new_n_n10_;
  assign new_n_n92_ = pv24_3_;
  assign pv119_17_ = new_n_n54_;
  assign pv151_20_ = new_n_n9_;
  assign new_n_n89_ = pv24_0_;
  assign new_n_n116_ = pv56_1_;
  assign pv119_14_ = new_n_n51_;
  assign pv151_23_ = new_n_n12_;
  assign new_n_n90_ = pv24_1_;
  assign new_n_n115_ = pv56_0_;
  assign new_n_n87_ = pv88_30_;
  assign pv119_15_ = new_n_n52_;
  assign pv151_22_ = new_n_n11_;
  assign new_n_n118_ = pv56_3_;
  assign new_n_n88_ = pv88_31_;
  assign pv119_12_ = new_n_n49_;
  assign pv151_25_ = new_n_n14_;
  assign pv151_30_ = new_n_n19_;
  assign new_n_n117_ = pv56_2_;
  assign pv119_13_ = new_n_n50_;
  assign pv151_24_ = new_n_n13_;
  assign pv151_31_ = new_n_n20_;
  assign new_n_n154_ = pv9_1_;
  assign new_n_n102_ = pv24_13_;
  assign pv119_10_ = new_n_n47_;
  assign pv151_5_ = new_n_n26_;
  assign pv151_14_ = new_n_n35_;
  assign new_n_n153_ = pv9_2_;
  assign new_n_n103_ = pv24_14_;
  assign pv119_11_ = new_n_n48_;
  assign pv151_4_ = new_n_n25_;
  assign pv151_15_ = new_n_n36_;
  assign new_n_n155_ = pv9_3_;
  assign new_n_n100_ = pv24_11_;
  assign new_n_n68_ = pv88_0_;
  assign pv151_7_ = new_n_n28_;
  assign pv151_12_ = new_n_n33_;
  assign new_n_n101_ = pv24_12_;
  assign new_n_n104_ = pv88_1_;
  assign pv151_6_ = new_n_n27_;
  assign pv151_13_ = new_n_n34_;
  assign new_n_n131_ = pv56_16_;
  assign new_n_n142_ = pv56_27_;
  assign pv151_9_ = new_n_n30_;
  assign pv151_10_ = new_n_n31_;
  assign new_n_n132_ = pv56_17_;
  assign new_n_n141_ = pv56_26_;
  assign pv151_8_ = new_n_n29_;
  assign pv151_11_ = new_n_n32_;
  assign new_n_n133_ = pv56_18_;
  assign new_n_n144_ = pv56_29_;
  assign new_n_n151_ = pv9_0_;
  assign new_n_n134_ = pv56_19_;
  assign new_n_n143_ = pv56_28_;
  assign new_nv158_ = new_nv157_ & new_nv155_ & new_nv156_;
  assign new_n_n3_ = new_nv168_ | new_nv170_ | new_nv171_ | new_nv169_ | new_nv165_ | new_nv167_;
  assign new_n_n63_ = new_nv212_ | new_nv267_ | new_nv236_ | new_nv180_ | new_nv437_;
  assign new_nv197_ = new_n_n125_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n41_ = new_nv207_ | new_nv289_ | new_nv377_ | new_nv202_ | new_nv437_;
  assign new_nv210_ = new_n_n136_ & new_nv207_;
  assign new_nv221_ = new_n_n125_ & new_nv207_;
  assign new_nv232_ = new_n_n135_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv243_ = new_n_n124_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv265_ = new_n_n129_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n21_ = new_nv296_ | new_nv295_ | new_nv425_ | new_nv294_ | new_nv329_ | new_nv297_ | new_nv393_ | new_nv361_;
  assign new_n_n10_ = new_nv296_ | new_nv295_ | new_nv404_ | new_nv294_ | new_nv308_ | new_nv297_ | new_nv372_ | new_nv340_;
  assign new_nv303_ = new_n_n83_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv314_ = new_n_n72_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv325_ = new_n_n107_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv336_ = new_n_n74_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv154_ = new_n_n153_ & new_n_n152_;
  assign new_n_n2_ = new_nv161_ | new_nv158_ | new_nv169_ | new_nv170_ | new_nv163_ | new_nv171_ | new_nv162_;
  assign new_nv180_ = new_n_n142_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv192_ = new_n_n130_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv203_ = new_n_n119_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv209_ = new_n_n137_ & new_nv207_;
  assign new_nv222_ = new_n_n124_ & new_nv207_;
  assign new_nv231_ = new_n_n115_ & new_nv207_;
  assign new_nv244_ = new_n_n123_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv264_ = new_n_n130_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n20_ = new_nv296_ | new_nv295_ | new_nv394_ | new_nv294_ | new_nv298_ | new_nv297_ | new_nv362_ | new_nv330_;
  assign new_n_n11_ = new_nv296_ | new_nv295_ | new_nv403_ | new_nv294_ | new_nv307_ | new_nv297_ | new_nv371_ | new_nv339_;
  assign new_nv304_ = new_n_n82_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv313_ = new_n_n73_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv326_ = new_n_n106_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv335_ = new_n_n75_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv162_ = new_nv157_ & new_nv155_ & new_n_n148_;
  assign new_nv171_ = new_n_n152_ & new_nv166_ & new_nv159_;
  assign new_n_n64_ = new_nv211_ | new_nv266_ | new_nv235_ | new_nv179_ | new_nv437_;
  assign new_n_n51_ = new_nv224_ | new_nv279_ | new_nv248_ | new_nv192_ | new_nv437_;
  assign new_nv198_ = new_n_n124_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv208_ = new_n_n138_ & new_nv207_;
  assign new_nv223_ = new_n_n123_ & new_nv207_;
  assign new_nv234_ = new_n_n133_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv241_ = new_n_n126_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv263_ = new_n_n131_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv289_ = new_n_n93_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n30_ = new_nv296_ | new_nv295_ | new_nv416_ | new_nv294_ | new_nv320_ | new_nv297_ | new_nv384_ | new_nv352_;
  assign new_nv305_ = new_n_n81_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv316_ = new_n_n70_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv323_ = new_n_n109_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv334_ = new_n_n76_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv161_ = new_nv157_ & new_n_n154_ & new_nv156_ & new_nv159_ & new_nv160_;
  assign new_n_n4_ = new_nv163_ | new_nv161_ | new_nv167_ | new_nv165_ | new_nv169_ | new_nv168_ | new_nv171_ | new_nv162_ | new_nv153_ | new_nv158_ | new_nv152_ | new_nv170_ | new_nv154_;
  assign new_nv179_ = new_n_n143_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv193_ = new_n_n129_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n46_ = new_nv229_ | new_nv284_ | new_nv372_ | new_nv197_ | new_nv437_;
  assign new_nv202_ = new_n_n120_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv224_ = new_n_n122_ & new_nv207_;
  assign new_nv233_ = new_n_n134_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv242_ = new_n_n125_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv251_ = new_n_n116_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv290_ = new_n_n92_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n31_ = new_nv296_ | new_nv295_ | new_nv415_ | new_nv294_ | new_nv319_ | new_nv297_ | new_nv383_ | new_nv351_;
  assign new_nv306_ = new_n_n80_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv315_ = new_n_n71_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv324_ = new_n_n108_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv333_ = new_n_n77_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv165_ = new_nv157_ & new_n_n154_ & new_nv164_ & new_n_n153_;
  assign new_n_n61_ = new_nv214_ | new_nv269_ | new_nv238_ | new_nv182_ | new_nv437_;
  assign new_nv188_ = new_n_n134_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv225_ = new_n_n121_ & new_nv207_;
  assign new_nv236_ = new_n_n131_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv247_ = new_n_n120_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv269_ = new_n_n125_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv280_ = new_n_n102_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv307_ = new_n_n79_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv318_ = new_n_n114_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv329_ = new_n_n68_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv340_ = new_n_n70_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv441_ = ~new_n_n2_;
  assign new_nv163_ = new_nv157_ & new_n_n154_ & new_n_n147_;
  assign new_nv183_ = new_n_n139_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n56_ = new_nv219_ | new_nv274_ | new_nv243_ | new_nv187_ | new_nv437_;
  assign new_nv226_ = new_n_n120_ & new_nv207_;
  assign new_nv235_ = new_n_n132_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv268_ = new_n_n126_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv270_ = new_n_n124_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv279_ = new_n_n103_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv308_ = new_n_n78_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv317_ = new_n_n69_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv330_ = new_n_n80_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv339_ = new_n_n71_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv176_ = new_n_n146_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n62_ = new_nv213_ | new_nv268_ | new_nv237_ | new_nv181_ | new_nv437_;
  assign new_nv187_ = new_n_n135_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv227_ = new_n_n119_ & new_nv207_;
  assign new_nv245_ = new_n_n122_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv267_ = new_n_n127_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv309_ = new_n_n77_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv320_ = new_n_n112_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv327_ = new_n_n105_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv338_ = new_n_n72_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_n_n67_ = new_nv208_ | new_nv263_ | new_nv232_ | new_nv176_ | new_nv437_;
  assign new_nv181_ = new_n_n141_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv182_ = new_n_n140_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv237_ = new_n_n130_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv246_ = new_n_n121_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv266_ = new_n_n128_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv310_ = new_n_n76_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv319_ = new_n_n113_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv328_ = new_n_n104_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv337_ = new_n_n73_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_n_n59_ = new_nv216_ | new_nv271_ | new_nv240_ | new_nv184_ | new_nv437_;
  assign new_nv190_ = new_n_n132_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n48_ = new_nv227_ | new_nv282_ | new_nv251_ | new_nv195_ | new_nv437_;
  assign new_nv201_ = new_n_n121_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n37_ = new_nv207_ | new_nv293_ | new_nv381_ | new_nv206_ | new_nv437_;
  assign new_nv273_ = new_n_n121_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv284_ = new_n_n98_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n35_ = new_nv296_ | new_nv295_ | new_nv411_ | new_nv294_ | new_nv315_ | new_nv297_ | new_nv379_ | new_nv347_;
  assign new_n_n24_ = new_nv296_ | new_nv295_ | new_nv422_ | new_nv294_ | new_nv326_ | new_nv297_ | new_nv390_ | new_nv358_;
  assign new_n_n13_ = new_nv296_ | new_nv295_ | new_nv401_ | new_nv294_ | new_nv305_ | new_nv297_ | new_nv369_ | new_nv337_;
  assign new_nv300_ = new_n_n86_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv164_ = ~new_n_n155_;
  assign new_nv185_ = new_n_n137_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n54_ = new_nv221_ | new_nv276_ | new_nv245_ | new_nv189_ | new_nv437_;
  assign new_nv196_ = new_n_n126_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n43_ = new_nv207_ | new_nv287_ | new_nv375_ | new_nv200_ | new_nv437_;
  assign new_nv217_ = new_n_n129_ & new_nv207_;
  assign new_nv274_ = new_n_n120_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv283_ = new_n_n99_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n34_ = new_nv296_ | new_nv295_ | new_nv412_ | new_nv294_ | new_nv316_ | new_nv297_ | new_nv380_ | new_nv348_;
  assign new_n_n25_ = new_nv296_ | new_nv295_ | new_nv421_ | new_nv294_ | new_nv325_ | new_nv297_ | new_nv389_ | new_nv357_;
  assign new_n_n12_ = new_nv296_ | new_nv295_ | new_nv402_ | new_nv294_ | new_nv306_ | new_nv297_ | new_nv370_ | new_nv338_;
  assign new_nv299_ = new_n_n87_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv166_ = ~new_n_n154_;
  assign new_n_n60_ = new_nv215_ | new_nv270_ | new_nv239_ | new_nv183_ | new_nv437_;
  assign new_nv189_ = new_n_n133_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n47_ = new_nv228_ | new_nv283_ | new_nv371_ | new_nv196_ | new_nv437_;
  assign new_n_n38_ = new_nv207_ | new_nv292_ | new_nv380_ | new_nv205_ | new_nv437_;
  assign new_nv216_ = new_n_n130_ & new_nv207_;
  assign new_nv271_ = new_n_n123_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv282_ = new_n_n100_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n33_ = new_nv296_ | new_nv295_ | new_nv413_ | new_nv294_ | new_nv317_ | new_nv297_ | new_nv381_ | new_nv349_;
  assign new_n_n22_ = new_nv296_ | new_nv295_ | new_nv424_ | new_nv294_ | new_nv328_ | new_nv297_ | new_nv392_ | new_nv360_;
  assign new_n_n15_ = new_nv296_ | new_nv295_ | new_nv399_ | new_nv294_ | new_nv303_ | new_nv297_ | new_nv367_ | new_nv335_;
  assign new_nv298_ = new_n_n88_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv437_ = ~new_n_n4_;
  assign new_nv184_ = new_n_n138_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n55_ = new_nv220_ | new_nv275_ | new_nv244_ | new_nv188_ | new_nv437_;
  assign new_n_n42_ = new_nv207_ | new_nv288_ | new_nv376_ | new_nv201_ | new_nv437_;
  assign new_nv206_ = new_n_n116_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv215_ = new_n_n131_ & new_nv207_;
  assign new_nv272_ = new_n_n122_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv281_ = new_n_n101_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n32_ = new_nv296_ | new_nv295_ | new_nv414_ | new_nv294_ | new_nv318_ | new_nv297_ | new_nv382_ | new_nv350_;
  assign new_n_n23_ = new_nv296_ | new_nv295_ | new_nv423_ | new_nv294_ | new_nv327_ | new_nv297_ | new_nv391_ | new_nv359_;
  assign new_n_n14_ = new_nv296_ | new_nv295_ | new_nv400_ | new_nv294_ | new_nv304_ | new_nv297_ | new_nv368_ | new_nv336_;
  assign new_n_n5_ = new_nv296_ | new_nv295_ | new_nv409_ | new_nv294_ | new_nv313_ | new_nv297_ | new_nv377_ | new_nv345_;
  assign new_nv440_ = ~new_n_n3_;
  assign new_nv169_ = new_nv160_ & new_nv166_ & new_nv156_ & new_nv159_;
  assign new_n_n65_ = new_nv210_ | new_nv265_ | new_nv234_ | new_nv178_ | new_nv437_;
  assign new_n_n57_ = new_nv218_ | new_nv273_ | new_nv242_ | new_nv186_ | new_nv437_;
  assign new_n_n50_ = new_nv225_ | new_nv280_ | new_nv249_ | new_nv193_ | new_nv437_;
  assign new_nv199_ = new_n_n123_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n39_ = new_nv207_ | new_nv291_ | new_nv379_ | new_nv204_ | new_nv437_;
  assign new_nv214_ = new_n_n132_ & new_nv207_;
  assign new_nv228_ = new_n_n118_ & new_nv207_;
  assign new_nv239_ = new_n_n128_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv250_ = new_n_n117_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv277_ = new_n_n117_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv288_ = new_n_n94_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv291_ = new_n_n91_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n28_ = new_nv296_ | new_nv295_ | new_nv418_ | new_nv294_ | new_nv322_ | new_nv297_ | new_nv386_ | new_nv354_;
  assign new_n_n17_ = new_nv296_ | new_nv295_ | new_nv397_ | new_nv294_ | new_nv301_ | new_nv297_ | new_nv365_ | new_nv333_;
  assign new_n_n6_ = new_nv296_ | new_nv295_ | new_nv408_ | new_nv294_ | new_nv312_ | new_nv297_ | new_nv376_ | new_nv344_;
  assign new_nv321_ = new_n_n111_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv332_ = new_n_n78_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv156_ = ~new_n_n150_;
  assign new_nv170_ = new_n_n148_ & new_nv166_ & new_nv159_;
  assign new_nv178_ = new_n_n144_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n52_ = new_nv223_ | new_nv278_ | new_nv247_ | new_nv191_ | new_nv437_;
  assign new_nv194_ = new_n_n128_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n45_ = new_nv230_ | new_nv285_ | new_nv373_ | new_nv198_ | new_nv437_;
  assign new_nv205_ = new_n_n117_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv213_ = new_n_n133_ & new_nv207_;
  assign new_nv218_ = new_n_n128_ & new_nv207_;
  assign new_nv240_ = new_n_n127_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv249_ = new_n_n118_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv278_ = new_n_n116_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv287_ = new_n_n95_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv292_ = new_n_n90_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n29_ = new_nv296_ | new_nv295_ | new_nv417_ | new_nv294_ | new_nv321_ | new_nv297_ | new_nv385_ | new_nv353_;
  assign new_n_n16_ = new_nv296_ | new_nv295_ | new_nv398_ | new_nv294_ | new_nv302_ | new_nv297_ | new_nv366_ | new_nv334_;
  assign new_n_n7_ = new_nv296_ | new_nv295_ | new_nv407_ | new_nv294_ | new_nv311_ | new_nv297_ | new_nv375_ | new_nv343_;
  assign new_nv322_ = new_n_n110_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv331_ = new_n_n79_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv157_ = ~new_n_n152_;
  assign new_nv153_ = new_n_n154_ & new_n_n152_;
  assign new_nv167_ = new_nv160_ & new_nv157_ & new_nv166_ & new_nv156_ & new_n_n151_ & new_n_n153_;
  assign new_n_n66_ = new_nv209_ | new_nv264_ | new_nv233_ | new_nv177_ | new_nv437_;
  assign new_n_n58_ = new_nv217_ | new_nv272_ | new_nv241_ | new_nv185_ | new_nv437_;
  assign new_nv191_ = new_n_n131_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n49_ = new_nv226_ | new_nv281_ | new_nv250_ | new_nv194_ | new_nv437_;
  assign new_nv200_ = new_n_n122_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n40_ = new_nv207_ | new_nv290_ | new_nv378_ | new_nv203_ | new_nv437_;
  assign new_nv212_ = new_n_n134_ & new_nv207_;
  assign new_nv219_ = new_n_n127_ & new_nv207_;
  assign new_nv230_ = new_n_n116_ & new_nv207_;
  assign new_nv248_ = new_n_n119_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv275_ = new_n_n119_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv286_ = new_n_n96_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv293_ = new_n_n89_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n26_ = new_nv296_ | new_nv295_ | new_nv420_ | new_nv294_ | new_nv324_ | new_nv297_ | new_nv388_ | new_nv356_;
  assign new_n_n19_ = new_nv296_ | new_nv295_ | new_nv395_ | new_nv294_ | new_nv299_ | new_nv297_ | new_nv363_ | new_nv331_;
  assign new_n_n8_ = new_nv296_ | new_nv295_ | new_nv406_ | new_nv294_ | new_nv310_ | new_nv297_ | new_nv374_ | new_nv342_;
  assign new_nv301_ = new_n_n85_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv312_ = new_n_n74_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv159_ = ~new_n_n153_;
  assign new_nv152_ = new_n_n155_ & new_n_n154_ & new_n_n153_;
  assign new_nv168_ = new_nv157_ & new_nv166_ & new_n_n147_ & new_n_n153_;
  assign new_nv177_ = new_n_n145_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv186_ = new_n_n136_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n53_ = new_nv222_ | new_nv277_ | new_nv246_ | new_nv190_ | new_nv437_;
  assign new_nv195_ = new_n_n127_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_n_n44_ = new_nv231_ | new_nv286_ | new_nv374_ | new_nv199_ | new_nv437_;
  assign new_nv204_ = new_n_n118_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv211_ = new_n_n135_ & new_nv207_;
  assign new_nv220_ = new_n_n126_ & new_nv207_;
  assign new_nv229_ = new_n_n117_ & new_nv207_;
  assign new_nv238_ = new_n_n129_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv276_ = new_n_n118_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv285_ = new_n_n97_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_n_n36_ = new_nv296_ | new_nv295_ | new_nv410_ | new_nv294_ | new_nv314_ | new_nv297_ | new_nv378_ | new_nv346_;
  assign new_n_n27_ = new_nv296_ | new_nv295_ | new_nv419_ | new_nv294_ | new_nv323_ | new_nv297_ | new_nv387_ | new_nv355_;
  assign new_n_n18_ = new_nv296_ | new_nv295_ | new_nv396_ | new_nv294_ | new_nv300_ | new_nv297_ | new_nv364_ | new_nv332_;
  assign new_n_n9_ = new_nv296_ | new_nv295_ | new_nv405_ | new_nv294_ | new_nv309_ | new_nv297_ | new_nv373_ | new_nv341_;
  assign new_nv302_ = new_n_n84_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv311_ = new_n_n75_ & new_nv440_ & new_n_n4_ & new_nv441_;
  assign new_nv160_ = ~new_n_n149_;
  assign new_nv346_ = new_n_n110_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv357_ = new_n_n143_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv368_ = new_n_n71_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv379_ = new_n_n106_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv390_ = new_n_n139_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv345_ = new_n_n111_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv358_ = new_n_n142_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv367_ = new_n_n72_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv380_ = new_n_n105_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv389_ = new_n_n140_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv344_ = new_n_n112_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv359_ = new_n_n141_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv370_ = new_n_n69_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv377_ = new_n_n108_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv388_ = new_n_n141_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv343_ = new_n_n113_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv360_ = new_n_n140_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv369_ = new_n_n70_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv378_ = new_n_n107_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv387_ = new_n_n142_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv155_ = ~new_n_n151_;
  assign new_nv342_ = new_n_n114_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv397_ = new_n_n70_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv408_ = new_n_n105_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv419_ = new_n_n138_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv297_ = new_nv437_ & new_n_n3_ & new_n_n2_;
  assign new_nv341_ = new_n_n69_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv398_ = new_n_n69_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv407_ = new_n_n106_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv420_ = new_n_n137_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv296_ = new_nv437_ & new_n_n3_ & new_nv441_;
  assign new_nv399_ = new_n_n114_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv410_ = new_n_n68_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv417_ = new_n_n140_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv295_ = new_nv437_ & new_nv440_ & new_n_n2_;
  assign new_nv400_ = new_n_n113_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv409_ = new_n_n104_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv418_ = new_n_n139_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv294_ = new_nv437_ & new_nv440_ & new_nv441_;
  assign new_nv371_ = new_n_n114_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv382_ = new_n_n68_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv393_ = new_n_n136_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv404_ = new_n_n109_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv415_ = new_n_n142_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv207_ = new_n_n4_ & new_nv440_ & new_n_n2_;
  assign new_nv372_ = new_n_n113_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv381_ = new_n_n104_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv394_ = new_n_n73_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv403_ = new_n_n110_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv416_ = new_n_n141_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv425_ = new_n_n132_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv351_ = new_n_n105_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv362_ = new_n_n77_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv395_ = new_n_n72_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv406_ = new_n_n107_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv413_ = new_n_n144_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv424_ = new_n_n133_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv352_ = new_n_n104_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv361_ = new_n_n139_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv396_ = new_n_n71_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv405_ = new_n_n108_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv414_ = new_n_n143_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv423_ = new_n_n134_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv350_ = new_n_n106_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv353_ = new_n_n68_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv364_ = new_n_n75_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv375_ = new_n_n110_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv386_ = new_n_n143_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv411_ = new_n_n146_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv422_ = new_n_n135_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv349_ = new_n_n107_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv354_ = new_n_n146_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv363_ = new_n_n76_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv376_ = new_n_n109_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv385_ = new_n_n144_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv412_ = new_n_n145_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv421_ = new_n_n136_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv348_ = new_n_n108_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv355_ = new_n_n145_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv366_ = new_n_n73_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv373_ = new_n_n112_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv384_ = new_n_n145_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv391_ = new_n_n138_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv402_ = new_n_n111_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
  assign new_nv347_ = new_n_n109_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv356_ = new_n_n144_ & new_nv440_ & new_n_n4_ & new_n_n2_;
  assign new_nv365_ = new_n_n74_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv374_ = new_n_n111_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv383_ = new_n_n146_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv392_ = new_n_n137_ & new_n_n3_ & new_n_n4_ & new_nv441_;
  assign new_nv401_ = new_n_n112_ & new_n_n3_ & new_n_n4_ & new_n_n2_;
endmodule


