// Benchmark "top" written by ABC on Sat Apr  1 09:44:31 2023

module top ( 
    pv96_30_, pv128_5_, pv160_1_, pv160_12_, pv160_25_, pv96_31_, pv128_6_,
    pv160_2_, pv160_11_, pv160_26_, pv96_10_, pv96_21_, pv128_3_,
    pv160_14_, pv160_27_, pv192_0_, pv96_11_, pv96_20_, pv128_4_, pv160_0_,
    pv160_13_, pv160_28_, pv128_1_, pv160_5_, pv160_29_, pv128_2_,
    pv128_19_, pv160_6_, pv199_4_, pv160_3_, pv160_10_, pv128_0_, pv160_4_,
    pv32_7_, pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv128_29_, pv192_19_,
    pv199_1_, pv32_6_, pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv192_18_,
    pv199_0_, pv32_5_, pv192_17_, pv192_31_, pv199_3_, pv32_4_, pv192_16_,
    pv192_30_, pv32_3_, pv64_4_, pv96_5_, pv128_9_, pv192_15_, pv192_20_,
    pv32_2_, pv64_5_, pv96_4_, pv192_14_, pv192_21_, pv32_1_, pv64_2_,
    pv96_7_, pv128_7_, pv192_13_, pv32_0_, pv64_3_, pv96_6_, pv128_8_,
    pv192_12_, pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_,
    pv128_21_, pv192_11_, pv192_24_, pv32_11_, pv32_20_, pv64_9_, pv64_18_,
    pv64_27_, pv96_0_, pv128_22_, pv192_10_, pv192_25_, pv32_12_, pv32_23_,
    pv32_30_, pv64_6_, pv64_15_, pv64_26_, pv96_3_, pv128_10_, pv128_23_,
    pv192_22_, pv32_13_, pv32_22_, pv32_31_, pv64_7_, pv64_16_, pv64_25_,
    pv96_2_, pv128_24_, pv128_31_, pv192_23_, pv32_14_, pv32_25_,
    pv128_25_, pv192_28_, pv32_15_, pv32_24_, pv128_26_, pv192_9_,
    pv192_29_, pv195_0_, pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv128_27_,
    pv192_26_, pv32_8_, pv32_17_, pv32_26_, pv64_29_, pv128_28_, pv192_27_,
    pv64_20_, pv64_31_, pv96_16_, pv96_27_, pv128_16_, pv160_9_, pv160_30_,
    pv192_6_, pv194_0_, pv64_10_, pv96_17_, pv96_26_, pv128_15_, pv160_19_,
    pv192_5_, pv96_18_, pv96_29_, pv128_18_, pv160_7_, pv192_8_, pv96_19_,
    pv96_28_, pv128_17_, pv160_8_, pv160_20_, pv192_7_, pv194_1_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv128_12_, pv128_30_, pv160_16_,
    pv160_21_, pv192_2_, pv64_14_, pv64_23_, pv96_13_, pv96_22_, pv128_11_,
    pv160_15_, pv160_22_, pv192_1_, pv64_11_, pv64_22_, pv96_14_, pv96_25_,
    pv128_14_, pv160_18_, pv160_23_, pv192_4_, pv64_12_, pv64_21_,
    pv64_30_, pv96_15_, pv96_24_, pv128_13_, pv128_20_, pv160_17_,
    pv160_24_, pv160_31_, pv192_3_,
    pv227_10_, pv227_23_, pv266_6_, pv227_0_, pv227_24_, pv227_21_,
    pv266_4_, pv227_22_, pv266_5_, pv227_27_, pv259_0_, pv227_25_,
    pv259_2_, pv227_26_, pv259_1_, pv227_7_, pv227_18_, pv259_17_,
    pv227_8_, pv227_17_, pv259_16_, pv227_5_, pv227_16_, pv259_19_,
    pv227_6_, pv227_15_, pv259_18_, pv227_3_, pv227_14_, pv259_26_,
    pv266_2_, pv227_4_, pv227_13_, pv227_20_, pv259_27_, pv266_3_,
    pv227_1_, pv227_12_, pv259_28_, pv266_0_, pv227_2_, pv227_11_,
    pv259_29_, pv266_1_, pv259_22_, pv259_23_, pv259_11_, pv259_24_,
    pv259_10_, pv259_25_, pv259_13_, pv259_31_, pv259_12_, pv259_30_,
    pv227_9_, pv259_15_, pv259_20_, pv227_19_, pv259_14_, pv259_21_,
    pv259_4_, pv259_3_, pv259_6_, pv259_5_, pv259_8_, pv259_7_, pv259_9_  );
  input  pv96_30_, pv128_5_, pv160_1_, pv160_12_, pv160_25_, pv96_31_,
    pv128_6_, pv160_2_, pv160_11_, pv160_26_, pv96_10_, pv96_21_, pv128_3_,
    pv160_14_, pv160_27_, pv192_0_, pv96_11_, pv96_20_, pv128_4_, pv160_0_,
    pv160_13_, pv160_28_, pv128_1_, pv160_5_, pv160_29_, pv128_2_,
    pv128_19_, pv160_6_, pv199_4_, pv160_3_, pv160_10_, pv128_0_, pv160_4_,
    pv32_7_, pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv128_29_, pv192_19_,
    pv199_1_, pv32_6_, pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv192_18_,
    pv199_0_, pv32_5_, pv192_17_, pv192_31_, pv199_3_, pv32_4_, pv192_16_,
    pv192_30_, pv32_3_, pv64_4_, pv96_5_, pv128_9_, pv192_15_, pv192_20_,
    pv32_2_, pv64_5_, pv96_4_, pv192_14_, pv192_21_, pv32_1_, pv64_2_,
    pv96_7_, pv128_7_, pv192_13_, pv32_0_, pv64_3_, pv96_6_, pv128_8_,
    pv192_12_, pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_,
    pv128_21_, pv192_11_, pv192_24_, pv32_11_, pv32_20_, pv64_9_, pv64_18_,
    pv64_27_, pv96_0_, pv128_22_, pv192_10_, pv192_25_, pv32_12_, pv32_23_,
    pv32_30_, pv64_6_, pv64_15_, pv64_26_, pv96_3_, pv128_10_, pv128_23_,
    pv192_22_, pv32_13_, pv32_22_, pv32_31_, pv64_7_, pv64_16_, pv64_25_,
    pv96_2_, pv128_24_, pv128_31_, pv192_23_, pv32_14_, pv32_25_,
    pv128_25_, pv192_28_, pv32_15_, pv32_24_, pv128_26_, pv192_9_,
    pv192_29_, pv195_0_, pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv128_27_,
    pv192_26_, pv32_8_, pv32_17_, pv32_26_, pv64_29_, pv128_28_, pv192_27_,
    pv64_20_, pv64_31_, pv96_16_, pv96_27_, pv128_16_, pv160_9_, pv160_30_,
    pv192_6_, pv194_0_, pv64_10_, pv96_17_, pv96_26_, pv128_15_, pv160_19_,
    pv192_5_, pv96_18_, pv96_29_, pv128_18_, pv160_7_, pv192_8_, pv96_19_,
    pv96_28_, pv128_17_, pv160_8_, pv160_20_, pv192_7_, pv194_1_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv128_12_, pv128_30_, pv160_16_,
    pv160_21_, pv192_2_, pv64_14_, pv64_23_, pv96_13_, pv96_22_, pv128_11_,
    pv160_15_, pv160_22_, pv192_1_, pv64_11_, pv64_22_, pv96_14_, pv96_25_,
    pv128_14_, pv160_18_, pv160_23_, pv192_4_, pv64_12_, pv64_21_,
    pv64_30_, pv96_15_, pv96_24_, pv128_13_, pv128_20_, pv160_17_,
    pv160_24_, pv160_31_, pv192_3_;
  output pv227_10_, pv227_23_, pv266_6_, pv227_0_, pv227_24_, pv227_21_,
    pv266_4_, pv227_22_, pv266_5_, pv227_27_, pv259_0_, pv227_25_,
    pv259_2_, pv227_26_, pv259_1_, pv227_7_, pv227_18_, pv259_17_,
    pv227_8_, pv227_17_, pv259_16_, pv227_5_, pv227_16_, pv259_19_,
    pv227_6_, pv227_15_, pv259_18_, pv227_3_, pv227_14_, pv259_26_,
    pv266_2_, pv227_4_, pv227_13_, pv227_20_, pv259_27_, pv266_3_,
    pv227_1_, pv227_12_, pv259_28_, pv266_0_, pv227_2_, pv227_11_,
    pv259_29_, pv266_1_, pv259_22_, pv259_23_, pv259_11_, pv259_24_,
    pv259_10_, pv259_25_, pv259_13_, pv259_31_, pv259_12_, pv259_30_,
    pv227_9_, pv259_15_, pv259_20_, pv227_19_, pv259_14_, pv259_21_,
    pv259_4_, pv259_3_, pv259_6_, pv259_5_, pv259_8_, pv259_7_, pv259_9_;
  wire new_n_n185_, new_n_n224_, new_n_n156_, new_n_n167_, new_n_n180_,
    new_n_n186_, new_n_n225_, new_n_n157_, new_n_n166_, new_n_n181_,
    new_n_n286_, new_n_n297_, new_n_n222_, new_n_n169_, new_n_n182_,
    new_n_n187_, new_n_n287_, new_n_n296_, new_n_n223_, new_n_n155_,
    new_n_n168_, new_n_n135_, new_n_n220_, new_n_n160_, new_n_n136_,
    new_n_n221_, new_n_n238_, new_n_n161_, new_n_n246_, new_n_n158_,
    new_n_n165_, new_n_n219_, new_n_n159_, new_n_n311_, new_n_n322_,
    new_n_n216_, new_n_n248_, new_n_n285_, new_n_n147_, new_n_n206_,
    new_n_n333_, new_n_n310_, new_n_n323_, new_n_n215_, new_n_n249_,
    new_n_n284_, new_n_n205_, new_n_n331_, new_n_n309_, new_n_n204_,
    new_n_n142_, new_n_n149_, new_n_n308_, new_n_n203_, new_n_n141_,
    new_n_n307_, new_n_n252_, new_n_n281_, new_n_n228_, new_n_n202_,
    new_n_n207_, new_n_n306_, new_n_n253_, new_n_n280_, new_n_n201_,
    new_n_n208_, new_n_n305_, new_n_n250_, new_n_n283_, new_n_n226_,
    new_n_n200_, new_n_n304_, new_n_n251_, new_n_n282_, new_n_n227_,
    new_n_n199_, new_n_n314_, new_n_n325_, new_n_n256_, new_n_n265_,
    new_n_n151_, new_n_n277_, new_n_n240_, new_n_n198_, new_n_n211_,
    new_n_n315_, new_n_n324_, new_n_n257_, new_n_n266_, new_n_n275_,
    new_n_n276_, new_n_n241_, new_n_n197_, new_n_n212_, new_n_n316_,
    new_n_n327_, new_n_n217_, new_n_n254_, new_n_n263_, new_n_n274_,
    new_n_n279_, new_n_n229_, new_n_n242_, new_n_n209_, new_n_n317_,
    new_n_n326_, new_n_n218_, new_n_n255_, new_n_n264_, new_n_n273_,
    new_n_n278_, new_n_n243_, new_n_n150_, new_n_n210_, new_n_n318_,
    new_n_n329_, new_n_n244_, new_n_n139_, new_n_n319_, new_n_n328_,
    new_n_n245_, new_n_n196_, new_n_n140_, new_n_n145_, new_n_n313_,
    new_n_n320_, new_n_n332_, new_n_n267_, new_n_n247_, new_n_n213_,
    new_n_n312_, new_n_n321_, new_n_n330_, new_n_n152_, new_n_n146_,
    new_n_n214_, new_n_n268_, new_n_n154_, new_n_n292_, new_n_n303_,
    new_n_n235_, new_n_n164_, new_n_n137_, new_n_n193_, new_n_n143_,
    new_n_n258_, new_n_n293_, new_n_n302_, new_n_n234_, new_n_n174_,
    new_n_n192_, new_n_n294_, new_n_n184_, new_n_n237_, new_n_n162_,
    new_n_n195_, new_n_n295_, new_n_n183_, new_n_n236_, new_n_n163_,
    new_n_n175_, new_n_n194_, new_n_n144_, new_n_n261_, new_n_n272_,
    new_n_n288_, new_n_n299_, new_n_n231_, new_n_n148_, new_n_n171_,
    new_n_n176_, new_n_n189_, new_n_n262_, new_n_n271_, new_n_n289_,
    new_n_n298_, new_n_n230_, new_n_n170_, new_n_n177_, new_n_n188_,
    new_n_n259_, new_n_n270_, new_n_n290_, new_n_n301_, new_n_n233_,
    new_n_n173_, new_n_n178_, new_n_n191_, new_n_n260_, new_n_n269_,
    new_n_n153_, new_n_n291_, new_n_n300_, new_n_n232_, new_n_n239_,
    new_n_n172_, new_n_n179_, new_n_n138_, new_n_n190_, new_nv268_,
    new_nv290_, new_n_n132_, new_nv305_, new_n_n121_, new_nv316_,
    new_n_n110_, new_nv329_, new_nv340_, new_nv401_, new_nv413_,
    new_nv424_, new_nv435_, new_nv445_, new_n_n99_, new_nv456_, new_nv481_,
    new_nv492_, new_nv503_, new_nv546_, new_nv557_, new_nv568_, new_nv291_,
    new_nv299_, new_n_n126_, new_nv310_, new_n_n115_, new_nv321_,
    new_nv330_, new_nv339_, new_nv391_, new_nv414_, new_nv423_, new_nv436_,
    new_n_n105_, new_nv451_, new_n_n94_, new_nv482_, new_nv491_,
    new_nv504_, new_nv545_, new_nv558_, new_nv567_, new_nv292_,
    new_n_n131_, new_nv304_, new_n_n122_, new_nv317_, new_n_n109_,
    new_nv327_, new_nv338_, new_nv392_, new_nv403_, new_nv422_, new_nv437_,
    new_nv446_, new_n_n100_, new_nv455_, new_nv468_, new_n_n76_,
    new_nv505_, new_nv548_, new_nv555_, new_nv566_, new_nv293_, new_nv300_,
    new_n_n127_, new_nv309_, new_n_n114_, new_nv322_, new_nv328_,
    new_nv337_, new_nv393_, new_nv402_, new_nv412_, new_nv438_,
    new_n_n104_, new_nv450_, new_n_n95_, new_n_n81_, new_nv473_,
    new_nv506_, new_nv547_, new_nv556_, new_nv565_, new_nv272_, new_nv283_,
    new_nv318_, new_n_n108_, new_nv344_, new_nv383_, new_nv439_,
    new_nv447_, new_n_n97_, new_nv458_, new_n_n86_, new_nv539_, new_nv550_,
    new_nv561_, new_nv574_, new_n_n7_, new_nv273_, new_nv282_, new_n_n113_,
    new_nv323_, new_nv345_, new_nv382_, new_nv440_, new_n_n103_,
    new_n_n92_, new_n_n91_, new_nv463_, new_nv540_, new_nv549_, new_nv562_,
    new_nv572_, new_nv270_, new_nv281_, new_nv331_, new_nv342_, new_nv381_,
    new_nv441_, new_n_n98_, new_nv457_, new_nv541_, new_nv552_, new_nv559_,
    new_nv570_, new_nv269_, new_nv271_, new_nv280_, new_nv332_, new_nv341_,
    new_nv343_, new_n_n102_, new_nv452_, new_n_n93_, new_nv542_,
    new_nv551_, new_nv560_, new_nv569_, new_nv276_, new_nv287_, new_nv298_,
    new_n_n128_, new_nv348_, new_nv387_, new_nv398_, new_nv410_,
    new_nv421_, new_nv460_, new_n_n84_, new_nv471_, new_nv478_, new_nv489_,
    new_nv500_, new_n_n3_, new_nv277_, new_nv286_, new_n_n133_, new_nv303_,
    new_nv349_, new_nv386_, new_nv399_, new_nv408_, new_nv431_, new_n_n89_,
    new_nv465_, new_n_n78_, new_nv477_, new_nv490_, new_nv499_, new_n_n4_,
    new_nv274_, new_nv285_, new_nv308_, new_n_n118_, new_nv346_,
    new_nv385_, new_nv400_, new_nv419_, new_nv430_, new_nv459_, new_n_n85_,
    new_nv472_, new_nv480_, new_nv487_, new_nv498_, new_n_n5_, new_nv275_,
    new_nv284_, new_n_n123_, new_nv313_, new_nv347_, new_nv384_,
    new_nv411_, new_nv420_, new_nv429_, new_n_n90_, new_nv464_, new_n_n77_,
    new_nv479_, new_nv488_, new_nv497_, new_n_n6_, new_nv294_, new_n_n130_,
    new_nv307_, new_n_n119_, new_nv314_, new_n_n112_, new_nv325_,
    new_nv336_, new_nv352_, new_nv394_, new_nv405_, new_nv417_, new_nv428_,
    new_nv443_, new_n_n101_, new_nv454_, new_nv462_, new_n_n82_,
    new_nv469_, new_n_n75_, new_nv485_, new_nv496_, new_nv553_, new_nv564_,
    new_nv573_, new_nv295_, new_nv301_, new_n_n124_, new_nv312_,
    new_n_n117_, new_nv319_, new_nv326_, new_nv335_, new_nv390_,
    new_nv395_, new_nv404_, new_nv418_, new_nv427_, new_nv432_, new_nv449_,
    new_n_n96_, new_n_n87_, new_nv467_, new_n_n80_, new_nv474_, new_nv486_,
    new_nv495_, new_nv554_, new_nv563_, new_nv578_, new_nv278_, new_nv289_,
    new_nv297_, new_n_n129_, new_nv306_, new_n_n120_, new_nv315_,
    new_n_n111_, new_nv324_, new_nv334_, new_nv350_, new_nv389_,
    new_nv396_, new_nv407_, new_nv415_, new_nv426_, new_nv433_, new_nv444_,
    new_nv453_, new_nv461_, new_n_n83_, new_nv470_, new_nv476_, new_nv483_,
    new_nv494_, new_nv501_, new_nv544_, new_nv604_, new_nv279_, new_nv288_,
    new_n_n134_, new_nv302_, new_n_n125_, new_nv311_, new_n_n116_,
    new_nv320_, new_n_n107_, new_nv333_, new_nv351_, new_nv388_,
    new_nv397_, new_nv406_, new_nv416_, new_nv425_, new_nv434_,
    new_n_n106_, new_nv448_, new_n_n88_, new_nv466_, new_n_n79_,
    new_nv475_, new_nv484_, new_nv493_, new_nv502_, new_nv543_, new_n_n2_,
    new_nv580_, new_n_n68_, new_nv602_, new_n_n59_, new_n_n48_, new_n_n74_,
    new_nv586_, new_nv601_, new_n_n58_, new_n_n49_, new_nv579_, new_nv587_,
    new_nv605_, new_n_n61_, new_n_n50_, new_nv577_, new_nv588_, new_nv603_,
    new_n_n60_, new_n_n51_, new_nv571_, new_nv576_, new_n_n41_, new_n_n30_,
    new_n_n19_, new_n_n8_, new_nv575_, new_n_n40_, new_n_n31_, new_n_n18_,
    new_n_n9_, new_n_n39_, new_n_n28_, new_n_n21_, new_n_n10_, new_n_n38_,
    new_n_n29_, new_n_n20_, new_n_n11_, new_n_n67_, new_n_n56_, new_n_n45_,
    new_n_n34_, new_n_n23_, new_n_n12_, new_n_n66_, new_n_n57_, new_n_n44_,
    new_n_n35_, new_n_n22_, new_n_n13_, new_n_n71_, new_nv590_, new_n_n43_,
    new_n_n32_, new_n_n25_, new_n_n14_, new_nv583_, new_nv589_, new_n_n42_,
    new_n_n33_, new_n_n24_, new_n_n15_, new_nv582_, new_n_n70_, new_nv598_,
    new_n_n63_, new_n_n52_, new_n_n27_, new_n_n16_, new_n_n72_, new_nv584_,
    new_nv597_, new_n_n62_, new_n_n53_, new_n_n26_, new_n_n17_, new_nv581_,
    new_n_n69_, new_nv600_, new_n_n65_, new_n_n54_, new_n_n47_, new_n_n36_,
    new_n_n73_, new_nv585_, new_nv599_, new_n_n64_, new_n_n55_, new_n_n46_,
    new_n_n37_;
  assign new_n_n185_ = pv96_30_;
  assign new_n_n224_ = pv128_5_;
  assign new_n_n156_ = pv160_1_;
  assign new_n_n167_ = pv160_12_;
  assign new_n_n180_ = pv160_25_;
  assign pv227_10_ = new_n_n117_;
  assign pv227_23_ = new_n_n130_;
  assign pv266_6_ = new_n_n74_;
  assign new_n_n186_ = pv96_31_;
  assign new_n_n225_ = pv128_6_;
  assign new_n_n157_ = pv160_2_;
  assign new_n_n166_ = pv160_11_;
  assign new_n_n181_ = pv160_26_;
  assign pv227_0_ = new_n_n107_;
  assign pv227_24_ = new_n_n131_;
  assign new_n_n286_ = pv96_10_;
  assign new_n_n297_ = pv96_21_;
  assign new_n_n222_ = pv128_3_;
  assign new_n_n169_ = pv160_14_;
  assign new_n_n182_ = pv160_27_;
  assign new_n_n187_ = pv192_0_;
  assign pv227_21_ = new_n_n128_;
  assign pv266_4_ = new_n_n72_;
  assign new_n_n287_ = pv96_11_;
  assign new_n_n296_ = pv96_20_;
  assign new_n_n223_ = pv128_4_;
  assign new_n_n155_ = pv160_0_;
  assign new_n_n168_ = pv160_13_;
  assign new_n_n135_ = pv160_28_;
  assign pv227_22_ = new_n_n129_;
  assign pv266_5_ = new_n_n73_;
  assign new_n_n220_ = pv128_1_;
  assign new_n_n160_ = pv160_5_;
  assign new_n_n136_ = pv160_29_;
  assign pv227_27_ = new_n_n134_;
  assign pv259_0_ = new_n_n75_;
  assign new_n_n221_ = pv128_2_;
  assign new_n_n238_ = pv128_19_;
  assign new_n_n161_ = pv160_6_;
  assign new_n_n246_ = pv199_4_;
  assign new_n_n158_ = pv160_3_;
  assign new_n_n165_ = pv160_10_;
  assign pv227_25_ = new_n_n132_;
  assign pv259_2_ = new_n_n77_;
  assign new_n_n219_ = pv128_0_;
  assign new_n_n159_ = pv160_4_;
  assign pv227_26_ = new_n_n133_;
  assign pv259_1_ = new_n_n76_;
  assign new_n_n311_ = pv32_7_;
  assign new_n_n322_ = pv32_18_;
  assign new_n_n216_ = pv32_29_;
  assign new_n_n248_ = pv64_0_;
  assign new_n_n285_ = pv96_9_;
  assign new_n_n147_ = pv128_29_;
  assign new_n_n206_ = pv192_19_;
  assign new_n_n333_ = pv199_1_;
  assign pv227_7_ = new_n_n114_;
  assign pv227_18_ = new_n_n125_;
  assign pv259_17_ = new_n_n92_;
  assign new_n_n310_ = pv32_6_;
  assign new_n_n323_ = pv32_19_;
  assign new_n_n215_ = pv32_28_;
  assign new_n_n249_ = pv64_1_;
  assign new_n_n284_ = pv96_8_;
  assign new_n_n205_ = pv192_18_;
  assign new_n_n331_ = pv199_0_;
  assign pv227_8_ = new_n_n115_;
  assign pv227_17_ = new_n_n124_;
  assign pv259_16_ = new_n_n91_;
  assign new_n_n309_ = pv32_5_;
  assign new_n_n204_ = pv192_17_;
  assign new_n_n142_ = pv192_31_;
  assign new_n_n149_ = pv199_3_;
  assign pv227_5_ = new_n_n112_;
  assign pv227_16_ = new_n_n123_;
  assign pv259_19_ = new_n_n94_;
  assign new_n_n308_ = pv32_4_;
  assign new_n_n203_ = pv192_16_;
  assign new_n_n141_ = pv192_30_;
  assign pv227_6_ = new_n_n113_;
  assign pv227_15_ = new_n_n122_;
  assign pv259_18_ = new_n_n93_;
  assign new_n_n307_ = pv32_3_;
  assign new_n_n252_ = pv64_4_;
  assign new_n_n281_ = pv96_5_;
  assign new_n_n228_ = pv128_9_;
  assign new_n_n202_ = pv192_15_;
  assign new_n_n207_ = pv192_20_;
  assign pv227_3_ = new_n_n110_;
  assign pv227_14_ = new_n_n121_;
  assign pv259_26_ = new_n_n101_;
  assign pv266_2_ = new_n_n70_;
  assign new_n_n306_ = pv32_2_;
  assign new_n_n253_ = pv64_5_;
  assign new_n_n280_ = pv96_4_;
  assign new_n_n201_ = pv192_14_;
  assign new_n_n208_ = pv192_21_;
  assign pv227_4_ = new_n_n111_;
  assign pv227_13_ = new_n_n120_;
  assign pv227_20_ = new_n_n127_;
  assign pv259_27_ = new_n_n102_;
  assign pv266_3_ = new_n_n71_;
  assign new_n_n305_ = pv32_1_;
  assign new_n_n250_ = pv64_2_;
  assign new_n_n283_ = pv96_7_;
  assign new_n_n226_ = pv128_7_;
  assign new_n_n200_ = pv192_13_;
  assign pv227_1_ = new_n_n108_;
  assign pv227_12_ = new_n_n119_;
  assign pv259_28_ = new_n_n103_;
  assign pv266_0_ = new_n_n68_;
  assign new_n_n304_ = pv32_0_;
  assign new_n_n251_ = pv64_3_;
  assign new_n_n282_ = pv96_6_;
  assign new_n_n227_ = pv128_8_;
  assign new_n_n199_ = pv192_12_;
  assign pv227_2_ = new_n_n109_;
  assign pv227_11_ = new_n_n118_;
  assign pv259_29_ = new_n_n104_;
  assign pv266_1_ = new_n_n69_;
  assign new_n_n314_ = pv32_10_;
  assign new_n_n325_ = pv32_21_;
  assign new_n_n256_ = pv64_8_;
  assign new_n_n265_ = pv64_17_;
  assign new_n_n151_ = pv64_28_;
  assign new_n_n277_ = pv96_1_;
  assign new_n_n240_ = pv128_21_;
  assign new_n_n198_ = pv192_11_;
  assign new_n_n211_ = pv192_24_;
  assign pv259_22_ = new_n_n97_;
  assign new_n_n315_ = pv32_11_;
  assign new_n_n324_ = pv32_20_;
  assign new_n_n257_ = pv64_9_;
  assign new_n_n266_ = pv64_18_;
  assign new_n_n275_ = pv64_27_;
  assign new_n_n276_ = pv96_0_;
  assign new_n_n241_ = pv128_22_;
  assign new_n_n197_ = pv192_10_;
  assign new_n_n212_ = pv192_25_;
  assign pv259_23_ = new_n_n98_;
  assign new_n_n316_ = pv32_12_;
  assign new_n_n327_ = pv32_23_;
  assign new_n_n217_ = pv32_30_;
  assign new_n_n254_ = pv64_6_;
  assign new_n_n263_ = pv64_15_;
  assign new_n_n274_ = pv64_26_;
  assign new_n_n279_ = pv96_3_;
  assign new_n_n229_ = pv128_10_;
  assign new_n_n242_ = pv128_23_;
  assign new_n_n209_ = pv192_22_;
  assign pv259_11_ = new_n_n86_;
  assign pv259_24_ = new_n_n99_;
  assign new_n_n317_ = pv32_13_;
  assign new_n_n326_ = pv32_22_;
  assign new_n_n218_ = pv32_31_;
  assign new_n_n255_ = pv64_7_;
  assign new_n_n264_ = pv64_16_;
  assign new_n_n273_ = pv64_25_;
  assign new_n_n278_ = pv96_2_;
  assign new_n_n243_ = pv128_24_;
  assign new_n_n150_ = pv128_31_;
  assign new_n_n210_ = pv192_23_;
  assign pv259_10_ = new_n_n85_;
  assign pv259_25_ = new_n_n100_;
  assign new_n_n318_ = pv32_14_;
  assign new_n_n329_ = pv32_25_;
  assign new_n_n244_ = pv128_25_;
  assign new_n_n139_ = pv192_28_;
  assign pv259_13_ = new_n_n88_;
  assign pv259_31_ = new_n_n106_;
  assign new_n_n319_ = pv32_15_;
  assign new_n_n328_ = pv32_24_;
  assign new_n_n245_ = pv128_26_;
  assign new_n_n196_ = pv192_9_;
  assign new_n_n140_ = pv192_29_;
  assign new_n_n145_ = pv195_0_;
  assign pv259_12_ = new_n_n87_;
  assign pv259_30_ = new_n_n105_;
  assign new_n_n313_ = pv32_9_;
  assign new_n_n320_ = pv32_16_;
  assign new_n_n332_ = pv32_27_;
  assign new_n_n267_ = pv64_19_;
  assign new_n_n247_ = pv128_27_;
  assign new_n_n213_ = pv192_26_;
  assign pv227_9_ = new_n_n116_;
  assign pv259_15_ = new_n_n90_;
  assign pv259_20_ = new_n_n95_;
  assign new_n_n312_ = pv32_8_;
  assign new_n_n321_ = pv32_17_;
  assign new_n_n330_ = pv32_26_;
  assign new_n_n152_ = pv64_29_;
  assign new_n_n146_ = pv128_28_;
  assign new_n_n214_ = pv192_27_;
  assign pv227_19_ = new_n_n126_;
  assign pv259_14_ = new_n_n89_;
  assign pv259_21_ = new_n_n96_;
  assign new_n_n268_ = pv64_20_;
  assign new_n_n154_ = pv64_31_;
  assign new_n_n292_ = pv96_16_;
  assign new_n_n303_ = pv96_27_;
  assign new_n_n235_ = pv128_16_;
  assign new_n_n164_ = pv160_9_;
  assign new_n_n137_ = pv160_30_;
  assign new_n_n193_ = pv192_6_;
  assign new_n_n143_ = pv194_0_;
  assign pv259_4_ = new_n_n79_;
  assign new_n_n258_ = pv64_10_;
  assign new_n_n293_ = pv96_17_;
  assign new_n_n302_ = pv96_26_;
  assign new_n_n234_ = pv128_15_;
  assign new_n_n174_ = pv160_19_;
  assign new_n_n192_ = pv192_5_;
  assign pv259_3_ = new_n_n78_;
  assign new_n_n294_ = pv96_18_;
  assign new_n_n184_ = pv96_29_;
  assign new_n_n237_ = pv128_18_;
  assign new_n_n162_ = pv160_7_;
  assign new_n_n195_ = pv192_8_;
  assign pv259_6_ = new_n_n81_;
  assign new_n_n295_ = pv96_19_;
  assign new_n_n183_ = pv96_28_;
  assign new_n_n236_ = pv128_17_;
  assign new_n_n163_ = pv160_8_;
  assign new_n_n175_ = pv160_20_;
  assign new_n_n194_ = pv192_7_;
  assign new_n_n144_ = pv194_1_;
  assign pv259_5_ = new_n_n80_;
  assign new_n_n261_ = pv64_13_;
  assign new_n_n272_ = pv64_24_;
  assign new_n_n288_ = pv96_12_;
  assign new_n_n299_ = pv96_23_;
  assign new_n_n231_ = pv128_12_;
  assign new_n_n148_ = pv128_30_;
  assign new_n_n171_ = pv160_16_;
  assign new_n_n176_ = pv160_21_;
  assign new_n_n189_ = pv192_2_;
  assign pv259_8_ = new_n_n83_;
  assign new_n_n262_ = pv64_14_;
  assign new_n_n271_ = pv64_23_;
  assign new_n_n289_ = pv96_13_;
  assign new_n_n298_ = pv96_22_;
  assign new_n_n230_ = pv128_11_;
  assign new_n_n170_ = pv160_15_;
  assign new_n_n177_ = pv160_22_;
  assign new_n_n188_ = pv192_1_;
  assign pv259_7_ = new_n_n82_;
  assign new_n_n259_ = pv64_11_;
  assign new_n_n270_ = pv64_22_;
  assign new_n_n290_ = pv96_14_;
  assign new_n_n301_ = pv96_25_;
  assign new_n_n233_ = pv128_14_;
  assign new_n_n173_ = pv160_18_;
  assign new_n_n178_ = pv160_23_;
  assign new_n_n191_ = pv192_4_;
  assign new_n_n260_ = pv64_12_;
  assign new_n_n269_ = pv64_21_;
  assign new_n_n153_ = pv64_30_;
  assign new_n_n291_ = pv96_15_;
  assign new_n_n300_ = pv96_24_;
  assign new_n_n232_ = pv128_13_;
  assign new_n_n239_ = pv128_20_;
  assign new_n_n172_ = pv160_17_;
  assign new_n_n179_ = pv160_24_;
  assign new_n_n138_ = pv160_31_;
  assign new_n_n190_ = pv192_3_;
  assign pv259_9_ = new_n_n84_;
  assign new_nv268_ = new_n_n332_ & new_nv573_ & new_n_n331_;
  assign new_nv290_ = new_n_n309_ & new_nv573_ & new_n_n331_;
  assign new_n_n132_ = new_nv299_ | new_nv383_ | new_nv270_ | new_nv327_;
  assign new_nv305_ = new_n_n295_ & new_nv573_ & new_nv578_;
  assign new_n_n121_ = new_nv310_ | new_nv394_ | new_nv281_ | new_nv338_;
  assign new_nv316_ = new_n_n284_ & new_nv573_ & new_nv578_;
  assign new_n_n110_ = new_nv321_ | new_nv405_ | new_nv292_ | new_nv349_;
  assign new_nv329_ = new_n_n271_ & new_n_n333_ & new_n_n331_;
  assign new_nv340_ = new_n_n260_ & new_n_n333_ & new_n_n331_;
  assign new_nv401_ = new_n_n9_ & new_n_n333_ & new_nv578_;
  assign new_nv413_ = new_n_n243_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv424_ = new_n_n232_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv435_ = new_n_n221_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv445_ = new_n_n212_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n99_ = new_nv482_ | new_nv572_ | new_nv546_ | new_nv450_ | new_nv417_;
  assign new_nv456_ = new_n_n201_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv481_ = new_n_n176_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv492_ = new_n_n165_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv503_ = new_n_n154_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv546_ = new_n_n54_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv557_ = new_n_n43_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv568_ = new_n_n32_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv291_ = new_n_n308_ & new_nv573_ & new_n_n331_;
  assign new_nv299_ = new_n_n301_ & new_nv573_ & new_nv578_;
  assign new_n_n126_ = new_nv305_ | new_nv389_ | new_nv276_ | new_nv333_;
  assign new_nv310_ = new_n_n290_ & new_nv573_ & new_nv578_;
  assign new_n_n115_ = new_nv316_ | new_nv400_ | new_nv287_ | new_nv344_;
  assign new_nv321_ = new_n_n279_ & new_nv573_ & new_nv578_;
  assign new_nv330_ = new_n_n270_ & new_n_n333_ & new_n_n331_;
  assign new_nv339_ = new_n_n261_ & new_n_n333_ & new_n_n331_;
  assign new_nv391_ = new_n_n19_ & new_n_n333_ & new_nv578_;
  assign new_nv414_ = new_n_n242_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv423_ = new_n_n233_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv436_ = new_n_n220_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_n_n105_ = new_nv476_ | new_nv572_ | new_nv540_ | new_nv444_ | new_nv411_;
  assign new_nv451_ = new_n_n206_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n94_ = new_nv487_ | new_nv572_ | new_nv551_ | new_nv455_ | new_nv422_;
  assign new_nv482_ = new_n_n175_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv491_ = new_n_n166_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv504_ = new_n_n153_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv545_ = new_n_n55_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv558_ = new_n_n42_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv567_ = new_n_n33_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv292_ = new_n_n307_ & new_nv573_ & new_n_n331_;
  assign new_n_n131_ = new_nv300_ | new_nv384_ | new_nv271_ | new_nv328_;
  assign new_nv304_ = new_n_n296_ & new_nv573_ & new_nv578_;
  assign new_n_n122_ = new_nv309_ | new_nv393_ | new_nv280_ | new_nv337_;
  assign new_nv317_ = new_n_n283_ & new_nv573_ & new_nv578_;
  assign new_n_n109_ = new_nv322_ | new_nv406_ | new_nv293_ | new_nv350_;
  assign new_nv327_ = new_n_n273_ & new_n_n333_ & new_n_n331_;
  assign new_nv338_ = new_n_n262_ & new_n_n333_ & new_n_n331_;
  assign new_nv392_ = new_n_n18_ & new_n_n333_ & new_nv578_;
  assign new_nv403_ = new_n_n7_ & new_n_n333_ & new_nv578_;
  assign new_nv422_ = new_n_n234_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv437_ = new_n_n219_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv446_ = new_n_n211_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n100_ = new_nv481_ | new_nv572_ | new_nv545_ | new_nv449_ | new_nv416_;
  assign new_nv455_ = new_n_n202_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv468_ = new_n_n189_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n76_ = new_nv505_ | new_nv572_ | new_nv569_ | new_nv473_ | new_nv440_;
  assign new_nv505_ = new_n_n152_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv548_ = new_n_n52_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv555_ = new_n_n45_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv566_ = new_n_n34_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv293_ = new_n_n306_ & new_nv573_ & new_n_n331_;
  assign new_nv300_ = new_n_n300_ & new_nv573_ & new_nv578_;
  assign new_n_n127_ = new_nv304_ | new_nv388_ | new_nv275_ | new_nv332_;
  assign new_nv309_ = new_n_n291_ & new_nv573_ & new_nv578_;
  assign new_n_n114_ = new_nv317_ | new_nv401_ | new_nv288_ | new_nv345_;
  assign new_nv322_ = new_n_n278_ & new_nv573_ & new_nv578_;
  assign new_nv328_ = new_n_n272_ & new_n_n333_ & new_n_n331_;
  assign new_nv337_ = new_n_n263_ & new_n_n333_ & new_n_n331_;
  assign new_nv393_ = new_n_n17_ & new_n_n333_ & new_nv578_;
  assign new_nv402_ = new_n_n8_ & new_n_n333_ & new_nv578_;
  assign new_nv412_ = new_n_n244_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv438_ = new_n_n218_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_n_n104_ = new_nv477_ | new_nv572_ | new_nv541_ | new_nv445_ | new_nv412_;
  assign new_nv450_ = new_n_n207_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n95_ = new_nv486_ | new_nv572_ | new_nv550_ | new_nv454_ | new_nv421_;
  assign new_n_n81_ = new_nv500_ | new_nv572_ | new_nv564_ | new_nv468_ | new_nv435_;
  assign new_nv473_ = new_n_n184_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv506_ = new_n_n151_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv547_ = new_n_n53_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv556_ = new_n_n44_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv565_ = new_n_n35_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv272_ = new_n_n327_ & new_nv573_ & new_n_n331_;
  assign new_nv283_ = new_n_n316_ & new_nv573_ & new_n_n331_;
  assign new_nv318_ = new_n_n282_ & new_nv573_ & new_nv578_;
  assign new_n_n108_ = new_nv323_ | new_nv407_ | new_nv294_ | new_nv351_;
  assign new_nv344_ = new_n_n256_ & new_n_n333_ & new_n_n331_;
  assign new_nv383_ = new_n_n27_ & new_n_n333_ & new_nv578_;
  assign new_nv439_ = new_n_n217_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv447_ = new_n_n210_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n97_ = new_nv484_ | new_nv572_ | new_nv548_ | new_nv452_ | new_nv419_;
  assign new_nv458_ = new_n_n199_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n86_ = new_nv495_ | new_nv572_ | new_nv559_ | new_nv463_ | new_nv430_;
  assign new_nv539_ = new_n_n61_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv550_ = new_n_n50_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv561_ = new_n_n39_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv574_ = new_n_n150_ & new_nv573_ & new_n_n149_ & new_n_n331_;
  assign new_n_n7_ = ~new_n_n281_;
  assign new_nv273_ = new_n_n326_ & new_nv573_ & new_n_n331_;
  assign new_nv282_ = new_n_n317_ & new_nv573_ & new_n_n331_;
  assign new_n_n113_ = new_nv318_ | new_nv402_ | new_nv289_ | new_nv346_;
  assign new_nv323_ = new_n_n277_ & new_nv573_ & new_nv578_;
  assign new_nv345_ = new_n_n255_ & new_n_n333_ & new_n_n331_;
  assign new_nv382_ = new_n_n28_ & new_n_n333_ & new_nv578_;
  assign new_nv440_ = new_n_n216_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_n_n103_ = new_nv478_ | new_nv572_ | new_nv542_ | new_nv446_ | new_nv413_;
  assign new_n_n92_ = new_nv489_ | new_nv572_ | new_nv553_ | new_nv457_ | new_nv424_;
  assign new_n_n91_ = new_nv490_ | new_nv572_ | new_nv554_ | new_nv458_ | new_nv425_;
  assign new_nv463_ = new_n_n194_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv540_ = new_n_n60_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv549_ = new_n_n51_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv562_ = new_n_n38_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv572_ = new_nv571_ & new_n_n333_;
  assign new_nv270_ = new_n_n329_ & new_nv573_ & new_n_n331_;
  assign new_nv281_ = new_n_n318_ & new_nv573_ & new_n_n331_;
  assign new_nv331_ = new_n_n269_ & new_n_n333_ & new_n_n331_;
  assign new_nv342_ = new_n_n258_ & new_n_n333_ & new_n_n331_;
  assign new_nv381_ = new_n_n29_ & new_n_n333_ & new_nv578_;
  assign new_nv441_ = new_n_n215_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_n_n98_ = new_nv483_ | new_nv572_ | new_nv547_ | new_nv451_ | new_nv418_;
  assign new_nv457_ = new_n_n200_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv541_ = new_n_n59_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv552_ = new_n_n48_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv559_ = new_n_n41_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv570_ = new_n_n30_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv269_ = new_n_n330_ & new_nv573_ & new_n_n331_;
  assign new_nv271_ = new_n_n328_ & new_nv573_ & new_n_n331_;
  assign new_nv280_ = new_n_n319_ & new_nv573_ & new_n_n331_;
  assign new_nv332_ = new_n_n268_ & new_n_n333_ & new_n_n331_;
  assign new_nv341_ = new_n_n259_ & new_n_n333_ & new_n_n331_;
  assign new_nv343_ = new_n_n257_ & new_n_n333_ & new_n_n331_;
  assign new_n_n102_ = new_nv479_ | new_nv572_ | new_nv543_ | new_nv447_ | new_nv414_;
  assign new_nv452_ = new_n_n205_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n93_ = new_nv488_ | new_nv572_ | new_nv552_ | new_nv456_ | new_nv423_;
  assign new_nv542_ = new_n_n58_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv551_ = new_n_n49_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv560_ = new_n_n40_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv569_ = new_n_n31_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv276_ = new_n_n323_ & new_nv573_ & new_n_n331_;
  assign new_nv287_ = new_n_n312_ & new_nv573_ & new_n_n331_;
  assign new_nv298_ = new_n_n302_ & new_nv573_ & new_nv578_;
  assign new_n_n128_ = new_nv303_ | new_nv387_ | new_nv274_ | new_nv331_;
  assign new_nv348_ = new_n_n252_ & new_n_n333_ & new_n_n331_;
  assign new_nv387_ = new_n_n23_ & new_n_n333_ & new_nv578_;
  assign new_nv398_ = new_n_n12_ & new_n_n333_ & new_nv578_;
  assign new_nv410_ = new_n_n247_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv421_ = new_n_n235_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv460_ = new_n_n197_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n84_ = new_nv497_ | new_nv572_ | new_nv561_ | new_nv465_ | new_nv432_;
  assign new_nv471_ = new_n_n186_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv478_ = new_n_n179_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv489_ = new_n_n168_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv500_ = new_n_n157_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_n_n3_ = ~new_n_n277_;
  assign new_nv277_ = new_n_n322_ & new_nv573_ & new_n_n331_;
  assign new_nv286_ = new_n_n313_ & new_nv573_ & new_n_n331_;
  assign new_n_n133_ = new_nv298_ | new_nv382_ | new_nv269_ | new_nv326_;
  assign new_nv303_ = new_n_n297_ & new_nv573_ & new_nv578_;
  assign new_nv349_ = new_n_n251_ & new_n_n333_ & new_n_n331_;
  assign new_nv386_ = new_n_n24_ & new_n_n333_ & new_nv578_;
  assign new_nv399_ = new_n_n11_ & new_n_n333_ & new_nv578_;
  assign new_nv408_ = new_n_n2_ & new_n_n333_ & new_nv578_;
  assign new_nv431_ = new_n_n225_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_n_n89_ = new_nv492_ | new_nv572_ | new_nv556_ | new_nv460_ | new_nv427_;
  assign new_nv465_ = new_n_n192_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n78_ = new_nv503_ | new_nv572_ | new_nv567_ | new_nv471_ | new_nv438_;
  assign new_nv477_ = new_n_n180_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv490_ = new_n_n167_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv499_ = new_n_n158_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_n_n4_ = ~new_n_n278_;
  assign new_nv274_ = new_n_n325_ & new_nv573_ & new_n_n331_;
  assign new_nv285_ = new_n_n314_ & new_nv573_ & new_n_n331_;
  assign new_nv308_ = new_n_n292_ & new_nv573_ & new_nv578_;
  assign new_n_n118_ = new_nv313_ | new_nv397_ | new_nv284_ | new_nv341_;
  assign new_nv346_ = new_n_n254_ & new_n_n333_ & new_n_n331_;
  assign new_nv385_ = new_n_n25_ & new_n_n333_ & new_nv578_;
  assign new_nv400_ = new_n_n10_ & new_n_n333_ & new_nv578_;
  assign new_nv419_ = new_n_n237_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv430_ = new_n_n226_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv459_ = new_n_n198_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n85_ = new_nv496_ | new_nv572_ | new_nv560_ | new_nv464_ | new_nv431_;
  assign new_nv472_ = new_n_n185_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv480_ = new_n_n177_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv487_ = new_n_n170_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv498_ = new_n_n159_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_n_n5_ = ~new_n_n279_;
  assign new_nv275_ = new_n_n324_ & new_nv573_ & new_n_n331_;
  assign new_nv284_ = new_n_n315_ & new_nv573_ & new_n_n331_;
  assign new_n_n123_ = new_nv308_ | new_nv392_ | new_nv279_ | new_nv336_;
  assign new_nv313_ = new_n_n287_ & new_nv573_ & new_nv578_;
  assign new_nv347_ = new_n_n253_ & new_n_n333_ & new_n_n331_;
  assign new_nv384_ = new_n_n26_ & new_n_n333_ & new_nv578_;
  assign new_nv411_ = new_n_n245_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv420_ = new_n_n236_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv429_ = new_n_n227_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_n_n90_ = new_nv491_ | new_nv572_ | new_nv555_ | new_nv459_ | new_nv426_;
  assign new_nv464_ = new_n_n193_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n77_ = new_nv504_ | new_nv572_ | new_nv568_ | new_nv472_ | new_nv439_;
  assign new_nv479_ = new_n_n178_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv488_ = new_n_n169_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv497_ = new_n_n160_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_n_n6_ = ~new_n_n280_;
  assign new_nv294_ = new_n_n305_ & new_nv573_ & new_n_n331_;
  assign new_n_n130_ = new_nv301_ | new_nv385_ | new_nv272_ | new_nv329_;
  assign new_nv307_ = new_n_n293_ & new_nv573_ & new_nv578_;
  assign new_n_n119_ = new_nv312_ | new_nv396_ | new_nv283_ | new_nv340_;
  assign new_nv314_ = new_n_n286_ & new_nv573_ & new_nv578_;
  assign new_n_n112_ = new_nv319_ | new_nv403_ | new_nv290_ | new_nv347_;
  assign new_nv325_ = new_n_n275_ & new_n_n333_ & new_n_n331_;
  assign new_nv336_ = new_n_n264_ & new_n_n333_ & new_n_n331_;
  assign new_nv352_ = new_n_n248_ & new_n_n333_ & new_n_n331_;
  assign new_nv394_ = new_n_n16_ & new_n_n333_ & new_nv578_;
  assign new_nv405_ = new_n_n5_ & new_n_n333_ & new_nv578_;
  assign new_nv417_ = new_n_n239_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv428_ = new_n_n228_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv443_ = new_n_n214_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n101_ = new_nv480_ | new_nv572_ | new_nv544_ | new_nv448_ | new_nv415_;
  assign new_nv454_ = new_n_n203_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv462_ = new_n_n195_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n82_ = new_nv499_ | new_nv572_ | new_nv563_ | new_nv467_ | new_nv434_;
  assign new_nv469_ = new_n_n188_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n75_ = new_nv506_ | new_nv572_ | new_nv570_ | new_nv474_ | new_nv441_;
  assign new_nv485_ = new_n_n172_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv496_ = new_n_n161_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv553_ = new_n_n47_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv564_ = new_n_n36_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv573_ = ~new_n_n333_;
  assign new_nv295_ = new_n_n304_ & new_nv573_ & new_n_n331_;
  assign new_nv301_ = new_n_n299_ & new_nv573_ & new_nv578_;
  assign new_n_n124_ = new_nv307_ | new_nv391_ | new_nv278_ | new_nv335_;
  assign new_nv312_ = new_n_n288_ & new_nv573_ & new_nv578_;
  assign new_n_n117_ = new_nv314_ | new_nv398_ | new_nv285_ | new_nv342_;
  assign new_nv319_ = new_n_n281_ & new_nv573_ & new_nv578_;
  assign new_nv326_ = new_n_n274_ & new_n_n333_ & new_n_n331_;
  assign new_nv335_ = new_n_n265_ & new_n_n333_ & new_n_n331_;
  assign new_nv390_ = new_n_n20_ & new_n_n333_ & new_nv578_;
  assign new_nv395_ = new_n_n15_ & new_n_n333_ & new_nv578_;
  assign new_nv404_ = new_n_n6_ & new_n_n333_ & new_nv578_;
  assign new_nv418_ = new_n_n238_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv427_ = new_n_n229_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv432_ = new_n_n224_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv449_ = new_n_n208_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n96_ = new_nv485_ | new_nv572_ | new_nv549_ | new_nv453_ | new_nv420_;
  assign new_n_n87_ = new_nv494_ | new_nv572_ | new_nv558_ | new_nv462_ | new_nv429_;
  assign new_nv467_ = new_n_n190_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n80_ = new_nv501_ | new_nv572_ | new_nv565_ | new_nv469_ | new_nv436_;
  assign new_nv474_ = new_n_n183_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv486_ = new_n_n171_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv495_ = new_n_n162_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv554_ = new_n_n46_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv563_ = new_n_n37_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv578_ = ~new_n_n331_;
  assign new_nv278_ = new_n_n321_ & new_nv573_ & new_n_n331_;
  assign new_nv289_ = new_n_n310_ & new_nv573_ & new_n_n331_;
  assign new_nv297_ = new_n_n303_ & new_nv573_ & new_nv578_;
  assign new_n_n129_ = new_nv302_ | new_nv386_ | new_nv273_ | new_nv330_;
  assign new_nv306_ = new_n_n294_ & new_nv573_ & new_nv578_;
  assign new_n_n120_ = new_nv311_ | new_nv395_ | new_nv282_ | new_nv339_;
  assign new_nv315_ = new_n_n285_ & new_nv573_ & new_nv578_;
  assign new_n_n111_ = new_nv320_ | new_nv404_ | new_nv291_ | new_nv348_;
  assign new_nv324_ = new_n_n276_ & new_nv573_ & new_nv578_;
  assign new_nv334_ = new_n_n266_ & new_n_n333_ & new_n_n331_;
  assign new_nv350_ = new_n_n250_ & new_n_n333_ & new_n_n331_;
  assign new_nv389_ = new_n_n21_ & new_n_n333_ & new_nv578_;
  assign new_nv396_ = new_n_n14_ & new_n_n333_ & new_nv578_;
  assign new_nv407_ = new_n_n3_ & new_n_n333_ & new_nv578_;
  assign new_nv415_ = new_n_n241_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv426_ = new_n_n230_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv433_ = new_n_n223_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv444_ = new_n_n213_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv453_ = new_n_n204_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv461_ = new_n_n196_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n83_ = new_nv498_ | new_nv572_ | new_nv562_ | new_nv466_ | new_nv433_;
  assign new_nv470_ = new_n_n187_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_nv476_ = new_n_n181_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv483_ = new_n_n174_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv494_ = new_n_n163_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv501_ = new_n_n156_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv544_ = new_n_n56_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_nv604_ = ~new_n_n149_;
  assign new_nv279_ = new_n_n320_ & new_nv573_ & new_n_n331_;
  assign new_nv288_ = new_n_n311_ & new_nv573_ & new_n_n331_;
  assign new_n_n134_ = new_nv297_ | new_nv381_ | new_nv268_ | new_nv325_;
  assign new_nv302_ = new_n_n298_ & new_nv573_ & new_nv578_;
  assign new_n_n125_ = new_nv306_ | new_nv390_ | new_nv277_ | new_nv334_;
  assign new_nv311_ = new_n_n289_ & new_nv573_ & new_nv578_;
  assign new_n_n116_ = new_nv315_ | new_nv399_ | new_nv286_ | new_nv343_;
  assign new_nv320_ = new_n_n280_ & new_nv573_ & new_nv578_;
  assign new_n_n107_ = new_nv324_ | new_nv408_ | new_nv295_ | new_nv352_;
  assign new_nv333_ = new_n_n267_ & new_n_n333_ & new_n_n331_;
  assign new_nv351_ = new_n_n249_ & new_n_n333_ & new_n_n331_;
  assign new_nv388_ = new_n_n22_ & new_n_n333_ & new_nv578_;
  assign new_nv397_ = new_n_n13_ & new_n_n333_ & new_nv578_;
  assign new_nv406_ = new_n_n4_ & new_n_n333_ & new_nv578_;
  assign new_nv416_ = new_n_n240_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv425_ = new_n_n231_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_nv434_ = new_n_n222_ & new_nv573_ & new_n_n246_ & new_n_n331_;
  assign new_n_n106_ = new_nv475_ | new_nv572_ | new_nv539_ | new_nv443_ | new_nv410_;
  assign new_nv448_ = new_n_n209_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n88_ = new_nv493_ | new_nv572_ | new_nv557_ | new_nv461_ | new_nv428_;
  assign new_nv466_ = new_n_n191_ & new_nv573_ & new_n_n246_ & new_nv578_;
  assign new_n_n79_ = new_nv502_ | new_nv572_ | new_nv566_ | new_nv470_ | new_nv437_;
  assign new_nv475_ = new_n_n182_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv484_ = new_n_n173_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv493_ = new_n_n164_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv502_ = new_n_n155_ & new_n_n333_ & new_n_n246_ & new_n_n331_;
  assign new_nv543_ = new_n_n57_ & new_n_n333_ & new_n_n246_ & new_nv578_;
  assign new_n_n2_ = ~new_n_n276_;
  assign new_nv580_ = new_n_n144_ & new_nv573_ & new_n_n149_ & new_nv578_;
  assign new_n_n68_ = new_nv590_ | new_nv605_ | new_nv603_ | new_nv585_ | new_nv577_;
  assign new_nv602_ = new_n_n63_ & new_n_n333_ & new_n_n149_ & new_nv578_;
  assign new_n_n59_ = ~new_n_n212_;
  assign new_n_n48_ = ~new_n_n201_;
  assign new_n_n74_ = new_nv597_ | new_nv579_;
  assign new_nv586_ = new_n_n149_ & new_n_n333_ & new_n_n331_;
  assign new_nv601_ = new_n_n64_ & new_n_n333_ & new_n_n149_ & new_nv578_;
  assign new_n_n58_ = ~new_n_n211_;
  assign new_n_n49_ = ~new_n_n202_;
  assign new_nv579_ = new_n_n145_ & new_nv573_ & new_n_n149_ & new_nv578_;
  assign new_nv587_ = new_n_n138_ & new_nv586_;
  assign new_nv605_ = new_nv604_ & new_n_n333_;
  assign new_n_n61_ = ~new_n_n214_;
  assign new_n_n50_ = ~new_n_n203_;
  assign new_nv577_ = new_n_n146_ & new_nv573_ & new_n_n149_ & new_n_n331_;
  assign new_nv588_ = new_n_n137_ & new_nv586_;
  assign new_nv603_ = new_n_n62_ & new_n_n333_ & new_n_n149_ & new_nv578_;
  assign new_n_n60_ = ~new_n_n213_;
  assign new_n_n51_ = ~new_n_n204_;
  assign new_nv571_ = ~new_n_n246_;
  assign new_nv576_ = new_n_n147_ & new_nv573_ & new_n_n149_ & new_n_n331_;
  assign new_n_n41_ = ~new_n_n194_;
  assign new_n_n30_ = ~new_n_n183_;
  assign new_n_n19_ = ~new_n_n293_;
  assign new_n_n8_ = ~new_n_n282_;
  assign new_nv575_ = new_n_n148_ & new_nv573_ & new_n_n149_ & new_n_n331_;
  assign new_n_n40_ = ~new_n_n193_;
  assign new_n_n31_ = ~new_n_n184_;
  assign new_n_n18_ = ~new_n_n292_;
  assign new_n_n9_ = ~new_n_n283_;
  assign new_n_n39_ = ~new_n_n192_;
  assign new_n_n28_ = ~new_n_n302_;
  assign new_n_n21_ = ~new_n_n295_;
  assign new_n_n10_ = ~new_n_n284_;
  assign new_n_n38_ = ~new_n_n191_;
  assign new_n_n29_ = ~new_n_n303_;
  assign new_n_n20_ = ~new_n_n294_;
  assign new_n_n11_ = ~new_n_n285_;
  assign new_n_n67_ = ~new_n_n144_;
  assign new_n_n56_ = ~new_n_n209_;
  assign new_n_n45_ = ~new_n_n198_;
  assign new_n_n34_ = ~new_n_n187_;
  assign new_n_n23_ = ~new_n_n297_;
  assign new_n_n12_ = ~new_n_n286_;
  assign new_n_n66_ = ~new_n_n143_;
  assign new_n_n57_ = ~new_n_n210_;
  assign new_n_n44_ = ~new_n_n197_;
  assign new_n_n35_ = ~new_n_n188_;
  assign new_n_n22_ = ~new_n_n296_;
  assign new_n_n13_ = ~new_n_n287_;
  assign new_n_n71_ = new_nv587_ | new_nv605_ | new_nv600_ | new_nv582_ | new_nv574_;
  assign new_nv590_ = new_n_n135_ & new_nv586_;
  assign new_n_n43_ = ~new_n_n196_;
  assign new_n_n32_ = ~new_n_n185_;
  assign new_n_n25_ = ~new_n_n299_;
  assign new_n_n14_ = ~new_n_n288_;
  assign new_nv583_ = new_n_n141_ & new_nv573_ & new_n_n149_ & new_nv578_;
  assign new_nv589_ = new_n_n136_ & new_nv586_;
  assign new_n_n42_ = ~new_n_n195_;
  assign new_n_n33_ = ~new_n_n186_;
  assign new_n_n24_ = ~new_n_n298_;
  assign new_n_n15_ = ~new_n_n289_;
  assign new_nv582_ = new_n_n142_ & new_nv573_ & new_n_n149_ & new_nv578_;
  assign new_n_n70_ = new_nv588_ | new_nv605_ | new_nv601_ | new_nv583_ | new_nv575_;
  assign new_nv598_ = new_n_n67_ & new_n_n333_ & new_n_n149_ & new_nv578_;
  assign new_n_n63_ = ~new_n_n140_;
  assign new_n_n52_ = ~new_n_n205_;
  assign new_n_n27_ = ~new_n_n301_;
  assign new_n_n16_ = ~new_n_n290_;
  assign new_n_n72_ = new_nv581_ | new_nv599_ | new_nv605_ | new_nv586_;
  assign new_nv584_ = new_n_n140_ & new_nv573_ & new_n_n149_ & new_nv578_;
  assign new_nv597_ = new_n_n145_ & new_n_n333_ & new_n_n149_ & new_nv578_;
  assign new_n_n62_ = ~new_n_n139_;
  assign new_n_n53_ = ~new_n_n206_;
  assign new_n_n26_ = ~new_n_n300_;
  assign new_n_n17_ = ~new_n_n291_;
  assign new_nv581_ = new_n_n143_ & new_nv573_ & new_n_n149_ & new_nv578_;
  assign new_n_n69_ = new_nv589_ | new_nv605_ | new_nv602_ | new_nv584_ | new_nv576_;
  assign new_nv600_ = new_n_n65_ & new_n_n333_ & new_n_n149_ & new_nv578_;
  assign new_n_n65_ = ~new_n_n142_;
  assign new_n_n54_ = ~new_n_n207_;
  assign new_n_n47_ = ~new_n_n200_;
  assign new_n_n36_ = ~new_n_n189_;
  assign new_n_n73_ = new_nv580_ | new_nv598_ | new_nv605_ | new_nv586_;
  assign new_nv585_ = new_n_n139_ & new_nv573_ & new_n_n149_ & new_nv578_;
  assign new_nv599_ = new_n_n66_ & new_n_n333_ & new_n_n149_ & new_nv578_;
  assign new_n_n64_ = ~new_n_n141_;
  assign new_n_n55_ = ~new_n_n208_;
  assign new_n_n46_ = ~new_n_n199_;
  assign new_n_n37_ = ~new_n_n190_;
endmodule


