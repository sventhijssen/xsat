// Benchmark "top" written by ABC on Fri Mar 31 12:10:15 2023

module top ( 
    pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0, px,
    pi0, py, pj0, pz, pk0, pl0, pm0, pa, pb, pc, pd, pe, pf, pg, ph, pi,
    pj, pk, pl, pm, pn, po,
    pn0, po0, pp0  );
  input  pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw,
    ph0, px, pi0, py, pj0, pz, pk0, pl0, pm0, pa, pb, pc, pd, pe, pf, pg,
    ph, pi, pj, pk, pl, pm, pn, po;
  output pn0, po0, pp0;
  wire new_na0_, new_nq_, new_nb0_, new_nr_, new_nc0_, new_ns_, new_nd0_,
    new_nt_, new_ne0_, new_nu_, new_nf0_, new_nv_, new_ng0_, new_nw_,
    new_nh0_, new_nx_, new_ni0_, new_ny_, new_nj0_, new_nz_, new_nk0_,
    new_nl0_, new_nm0_, new_na_, new_nb_, new_nc_, new_nd_, new_ne_,
    new_nf_, new_ng_, new_nh_, new_ni_, new_nj_, new_nk_, new_nl_, new_nm_,
    new_nn_, new_no_, new_n_n1017_, new_n_n1006_, new_n_n995_, new_n_n984_,
    new_n_n973_, new_n_n962_, new_n_n953_, new_n_n942_, new_n_n931_,
    new_n_n920_, new_n_n909_, new_n_n898_, new_n_n854_, new_n_n843_,
    new_n_n832_, new_n_n821_, new_n_n810_, new_n_n799_, new_n_n788_,
    new_n_n756_, new_n_n745_, new_n_n734_, new_n_n723_, new_n_n712_,
    new_n_n701_, new_n_n690_, new_n_n679_, new_n_n657_, new_n_n646_,
    new_n_n635_, new_n_n624_, new_n_n613_, new_n_n602_, new_n_n591_,
    new_n_n580_, new_n_n569_, new_n_n558_, new_n_n548_, new_n_n537_,
    new_n_n526_, new_n_n515_, new_n_n504_, new_n_n493_, new_n_n482_,
    new_n_n471_, new_n_n460_, new_n_n449_, new_n_n438_, new_n_n427_,
    new_n_n416_, new_n_n405_, new_n_n394_, new_n_n383_, new_n_n372_,
    new_n_n361_, new_n_n339_, new_n_n328_, new_n_n317_, new_n_n306_,
    new_n_n295_, new_n_n284_, new_n_n273_, new_n_n262_, new_n_n229_,
    new_n_n218_, new_n_n207_, new_n_n196_, new_n_n185_, new_n_n174_,
    new_n_n163_, new_n_n119_, new_n_n108_, new_n_n97_, new_n_n86_,
    new_n_n75_, new_n_n64_, new_n_n1016_, new_n_n1007_, new_n_n994_,
    new_n_n985_, new_n_n972_, new_n_n963_, new_n_n952_, new_n_n943_,
    new_n_n930_, new_n_n921_, new_n_n908_, new_n_n899_, new_n_n853_,
    new_n_n844_, new_n_n831_, new_n_n822_, new_n_n809_, new_n_n800_,
    new_n_n779_, new_n_n755_, new_n_n746_, new_n_n733_, new_n_n724_,
    new_n_n711_, new_n_n702_, new_n_n689_, new_n_n680_, new_n_n656_,
    new_n_n647_, new_n_n634_, new_n_n625_, new_n_n612_, new_n_n603_,
    new_n_n590_, new_n_n581_, new_n_n559_, new_n_n557_, new_n_n549_,
    new_n_n536_, new_n_n527_, new_n_n514_, new_n_n505_, new_n_n492_,
    new_n_n483_, new_n_n470_, new_n_n461_, new_n_n459_, new_n_n437_,
    new_n_n428_, new_n_n415_, new_n_n406_, new_n_n393_, new_n_n384_,
    new_n_n371_, new_n_n362_, new_n_n338_, new_n_n329_, new_n_n316_,
    new_n_n307_, new_n_n294_, new_n_n285_, new_n_n272_, new_n_n263_,
    new_n_n239_, new_n_n217_, new_n_n208_, new_n_n195_, new_n_n186_,
    new_n_n173_, new_n_n164_, new_n_n118_, new_n_n109_, new_n_n96_,
    new_n_n87_, new_n_n74_, new_n_n65_, new_n_n1026_, new_n_n993_,
    new_n_n982_, new_n_n975_, new_n_n964_, new_n_n955_, new_n_n944_,
    new_n_n929_, new_n_n918_, new_n_n911_, new_n_n900_, new_n_n856_,
    new_n_n845_, new_n_n830_, new_n_n819_, new_n_n812_, new_n_n801_,
    new_n_n769_, new_n_n758_, new_n_n747_, new_n_n732_, new_n_n721_,
    new_n_n714_, new_n_n703_, new_n_n670_, new_n_n659_, new_n_n648_,
    new_n_n633_, new_n_n622_, new_n_n615_, new_n_n604_, new_n_n589_,
    new_n_n571_, new_n_n560_, new_n_n535_, new_n_n524_, new_n_n517_,
    new_n_n506_, new_n_n491_, new_n_n480_, new_n_n473_, new_n_n462_,
    new_n_n436_, new_n_n425_, new_n_n418_, new_n_n407_, new_n_n392_,
    new_n_n381_, new_n_n374_, new_n_n363_, new_n_n337_, new_n_n326_,
    new_n_n319_, new_n_n308_, new_n_n293_, new_n_n282_, new_n_n275_,
    new_n_n264_, new_n_n238_, new_n_n227_, new_n_n209_, new_n_n194_,
    new_n_n183_, new_n_n176_, new_n_n165_, new_n_n139_, new_n_n128_,
    new_n_n95_, new_n_n84_, new_n_n77_, new_n_n66_, new_n_n1027_,
    new_n_n992_, new_n_n983_, new_n_n974_, new_n_n965_, new_n_n954_,
    new_n_n945_, new_n_n928_, new_n_n919_, new_n_n910_, new_n_n901_,
    new_n_n855_, new_n_n846_, new_n_n829_, new_n_n820_, new_n_n811_,
    new_n_n802_, new_n_n759_, new_n_n757_, new_n_n748_, new_n_n731_,
    new_n_n722_, new_n_n713_, new_n_n704_, new_n_n669_, new_n_n660_,
    new_n_n658_, new_n_n632_, new_n_n623_, new_n_n614_, new_n_n605_,
    new_n_n579_, new_n_n570_, new_n_n561_, new_n_n534_, new_n_n525_,
    new_n_n516_, new_n_n507_, new_n_n490_, new_n_n481_, new_n_n472_,
    new_n_n463_, new_n_n435_, new_n_n426_, new_n_n417_, new_n_n408_,
    new_n_n391_, new_n_n382_, new_n_n373_, new_n_n364_, new_n_n336_,
    new_n_n327_, new_n_n318_, new_n_n309_, new_n_n292_, new_n_n283_,
    new_n_n274_, new_n_n265_, new_n_n237_, new_n_n228_, new_n_n219_,
    new_n_n193_, new_n_n184_, new_n_n175_, new_n_n166_, new_n_n138_,
    new_n_n129_, new_n_n94_, new_n_n85_, new_n_n76_, new_n_n67_,
    new_n_n1024_, new_n_n1013_, new_n_n1002_, new_n_n977_, new_n_n966_,
    new_n_n949_, new_n_n938_, new_n_n935_, new_n_n924_, new_n_n913_,
    new_n_n902_, new_n_n850_, new_n_n839_, new_n_n836_, new_n_n825_,
    new_n_n814_, new_n_n803_, new_n_n752_, new_n_n741_, new_n_n738_,
    new_n_n727_, new_n_n716_, new_n_n705_, new_n_n653_, new_n_n642_,
    new_n_n628_, new_n_n617_, new_n_n606_, new_n_n554_, new_n_n544_,
    new_n_n519_, new_n_n508_, new_n_n456_, new_n_n445_, new_n_n409_,
    new_n_n390_, new_n_n357_, new_n_n346_, new_n_n291_, new_n_n280_,
    new_n_n258_, new_n_n247_, new_n_n192_, new_n_n181_, new_n_n170_,
    new_n_n159_, new_n_n148_, new_n_n93_, new_n_n82_, new_n_n71_,
    new_n_n60_, new_n_n9_, new_n_n1025_, new_n_n1012_, new_n_n1003_,
    new_n_n976_, new_n_n967_, new_n_n948_, new_n_n939_, new_n_n934_,
    new_n_n925_, new_n_n912_, new_n_n903_, new_n_n849_, new_n_n840_,
    new_n_n835_, new_n_n826_, new_n_n813_, new_n_n804_, new_n_n751_,
    new_n_n742_, new_n_n737_, new_n_n728_, new_n_n715_, new_n_n706_,
    new_n_n652_, new_n_n643_, new_n_n638_, new_n_n616_, new_n_n607_,
    new_np0_, new_n_n545_, new_n_n518_, new_n_n509_, new_n_n455_,
    new_n_n446_, new_n_n419_, new_n_n380_, new_n_n356_, new_n_n347_,
    new_n_n290_, new_n_n281_, new_n_n257_, new_n_n248_, new_n_n191_,
    new_n_n182_, new_n_n160_, new_n_n158_, new_n_n149_, new_n_n92_,
    new_n_n83_, new_n_n70_, new_n_n61_, new_n_n1022_, new_n_n1015_,
    new_n_n1004_, new_n_n997_, new_n_n986_, new_n_n951_, new_n_n940_,
    new_n_n933_, new_n_n922_, new_n_n915_, new_n_n904_, new_n_n852_,
    new_n_n841_, new_n_n834_, new_n_n823_, new_n_n816_, new_n_n805_,
    new_n_n754_, new_n_n743_, new_n_n736_, new_n_n725_, new_n_n718_,
    new_n_n707_, new_n_n655_, new_n_n644_, new_n_n637_, new_n_n626_,
    new_n_n608_, new_n_n556_, new_n_n546_, new_n_n539_, new_n_n528_,
    new_n_n458_, new_n_n447_, new_n_n429_, new_n_n370_, new_n_n359_,
    new_n_n348_, new_n_n271_, new_n_n260_, new_n_n249_, new_n_n190_,
    new_n_n172_, new_n_n161_, new_n_n91_, new_n_n80_, new_n_n73_,
    new_n_n62_, new_n_n1023_, new_n_n1014_, new_n_n1005_, new_n_n996_,
    new_n_n987_, new_n_n950_, new_n_n941_, new_n_n932_, new_n_n923_,
    new_n_n914_, new_n_n905_, new_n_n851_, new_n_n842_, new_n_n833_,
    new_n_n824_, new_n_n815_, new_n_n806_, new_n_n753_, new_n_n744_,
    new_n_n735_, new_n_n726_, new_n_n717_, new_n_n708_, new_n_n654_,
    new_n_n645_, new_n_n636_, new_n_n627_, new_n_n618_, new_n_n555_,
    new_n_n547_, new_n_n538_, new_n_n529_, new_n_n457_, new_n_n448_,
    new_n_n439_, new_n_n360_, new_n_n358_, new_n_n349_, new_n_n270_,
    new_n_n261_, new_n_n259_, new_n_n180_, new_n_n171_, new_n_n162_,
    new_n_n90_, new_n_n81_, new_n_n72_, new_n_n63_, new_n_n895_,
    new_n_n884_, new_n_n873_, new_n_n862_, new_n_n796_, new_n_n786_,
    new_n_n775_, new_n_n764_, new_n_n698_, new_n_n687_, new_n_n676_,
    new_n_n665_, new_n_n649_, new_n_n588_, new_n_n577_, new_n_n566_,
    new_n_n551_, new_n_n540_, new_n_n479_, new_n_n468_, new_n_n452_,
    new_n_n441_, new_n_n430_, new_n_n369_, new_n_n353_, new_n_n342_,
    new_n_n331_, new_n_n320_, new_n_n254_, new_n_n243_, new_n_n232_,
    new_n_n221_, new_n_n210_, new_n_n155_, new_n_n144_, new_n_n133_,
    new_n_n122_, new_n_n111_, new_n_n100_, new_n_n5_, new_n_n894_,
    new_n_n885_, new_n_n872_, new_n_n863_, new_n_n795_, new_n_n787_,
    new_n_n774_, new_n_n765_, new_n_n697_, new_n_n688_, new_n_n675_,
    new_n_n666_, new_n_n639_, new_n_n598_, new_n_n576_, new_n_n567_,
    new_n_n550_, new_n_n541_, new_n_n478_, new_n_n469_, new_n_n451_,
    new_n_n442_, new_n_n420_, new_n_n379_, new_n_n352_, new_n_n343_,
    new_n_n330_, new_n_n321_, new_n_n253_, new_n_n244_, new_n_n231_,
    new_n_n222_, new_n_n200_, new_n_n154_, new_n_n145_, new_n_n132_,
    new_n_n123_, new_n_n110_, new_n_n101_, new_n_n6_, new_n_n893_,
    new_n_n882_, new_n_n875_, new_n_n864_, new_n_n848_, new_n_n794_,
    new_n_n784_, new_n_n777_, new_n_n766_, new_n_n750_, new_n_n739_,
    new_n_n696_, new_n_n685_, new_n_n678_, new_n_n667_, new_n_n651_,
    new_n_n640_, new_n_n597_, new_n_n586_, new_n_n568_, new_n_n553_,
    new_n_n542_, new_n_n499_, new_n_n488_, new_n_n454_, new_n_n443_,
    new_n_n410_, new_n_n389_, new_n_n355_, new_n_n344_, new_n_n311_,
    new_n_n300_, new_n_n256_, new_n_n245_, new_n_n230_, new_n_n212_,
    new_n_n201_, new_n_n157_, new_n_n146_, new_n_n131_, new_n_n120_,
    new_n_n113_, new_n_n102_, new_n_n7_, new_n_n892_, new_n_n883_,
    new_n_n874_, new_n_n865_, new_n_n838_, new_n_n793_, new_n_n785_,
    new_n_n776_, new_n_n767_, new_n_n749_, new_n_n740_, new_n_n695_,
    new_n_n686_, new_n_n677_, new_n_n668_, new_n_n650_, new_n_n641_,
    new_n_n596_, new_n_n587_, new_n_n578_, new_n_n552_, new_n_n543_,
    new_n_n498_, new_n_n489_, new_n_n453_, new_n_n444_, new_n_n400_,
    new_n_n399_, new_n_n354_, new_n_n345_, new_n_n310_, new_n_n301_,
    new_n_n255_, new_n_n246_, new_n_n220_, new_n_n211_, new_n_n202_,
    new_n_n156_, new_n_n147_, new_n_n130_, new_n_n121_, new_n_n112_,
    new_n_n103_, new_n_n8_, new_n_n891_, new_n_n880_, new_n_n869_,
    new_n_n858_, new_n_n828_, new_n_n792_, new_n_n782_, new_n_n771_,
    new_n_n760_, new_n_n730_, new_n_n719_, new_n_n694_, new_n_n683_,
    new_n_n672_, new_n_n661_, new_n_n631_, new_n_n620_, new_n_n609_,
    new_n_n595_, new_n_n584_, new_n_n573_, new_n_n562_, new_n_n533_,
    new_n_n522_, new_n_n511_, new_n_n500_, new_n_n497_, new_n_n486_,
    new_n_n475_, new_n_n464_, new_n_n434_, new_n_n423_, new_n_n412_,
    new_n_n401_, new_n_n398_, new_n_n387_, new_n_n376_, new_n_n365_,
    new_n_n335_, new_n_n324_, new_n_n313_, new_n_n302_, new_n_n299_,
    new_n_n288_, new_n_n277_, new_n_n266_, new_n_n250_, new_n_n236_,
    new_n_n225_, new_n_n214_, new_n_n203_, new_n_n189_, new_n_n178_,
    new_n_n167_, new_n_n151_, new_n_n140_, new_n_n137_, new_n_n126_,
    new_n_n115_, new_n_n104_, new_n_n79_, new_n_n68_, new_n_n1_,
    new_n_n890_, new_n_n881_, new_n_n868_, new_n_n859_, new_n_n818_,
    new_n_n791_, new_n_n783_, new_n_n770_, new_n_n761_, new_n_n729_,
    new_n_n720_, new_n_n693_, new_n_n684_, new_n_n671_, new_n_n662_,
    new_n_n630_, new_n_n621_, new_n_n599_, new_n_n594_, new_n_n585_,
    new_n_n572_, new_n_n563_, new_n_n532_, new_n_n523_, new_n_n510_,
    new_n_n501_, new_n_n496_, new_n_n487_, new_n_n474_, new_n_n465_,
    new_n_n433_, new_n_n424_, new_n_n411_, new_n_n402_, new_n_n397_,
    new_n_n388_, new_n_n375_, new_n_n366_, new_n_n334_, new_n_n325_,
    new_n_n312_, new_n_n303_, new_n_n298_, new_n_n289_, new_n_n276_,
    new_n_n267_, new_n_n240_, new_n_n235_, new_n_n226_, new_n_n213_,
    new_n_n204_, new_n_n199_, new_n_n177_, new_n_n168_, new_n_n150_,
    new_n_n141_, new_n_n136_, new_n_n127_, new_n_n114_, new_n_n105_,
    new_n_n78_, new_n_n69_, new_n_n2_, new_n_n889_, new_n_n878_,
    new_n_n871_, new_n_n860_, new_n_n808_, new_n_n790_, new_n_n780_,
    new_n_n773_, new_n_n762_, new_n_n710_, new_n_n699_, new_n_n692_,
    new_n_n681_, new_n_n674_, new_n_n663_, new_n_n629_, new_n_n611_,
    new_n_n600_, new_n_n593_, new_n_n582_, new_n_n575_, new_n_n564_,
    new_n_n531_, new_n_n520_, new_n_n513_, new_n_n502_, new_n_n495_,
    new_n_n484_, new_n_n477_, new_n_n466_, new_n_n450_, new_n_n432_,
    new_n_n421_, new_n_n414_, new_n_n403_, new_n_n396_, new_n_n385_,
    new_n_n378_, new_n_n367_, new_n_n351_, new_n_n340_, new_n_n333_,
    new_n_n322_, new_n_n315_, new_n_n304_, new_n_n297_, new_n_n286_,
    new_n_n279_, new_n_n268_, new_n_n252_, new_n_n241_, new_n_n234_,
    new_n_n223_, new_n_n216_, new_n_n205_, new_n_n198_, new_n_n187_,
    new_n_n169_, new_n_n153_, new_n_n142_, new_n_n135_, new_n_n124_,
    new_n_n117_, new_n_n106_, new_n_n99_, new_n_n88_, new_n_n3_,
    new_n_n888_, new_n_n879_, new_n_n870_, new_n_n861_, new_n_n798_,
    new_n_n789_, new_n_n781_, new_n_n772_, new_n_n763_, new_n_n709_,
    new_n_n700_, new_n_n691_, new_n_n682_, new_n_n673_, new_n_n664_,
    new_n_n619_, new_n_n610_, new_n_n601_, new_n_n592_, new_n_n583_,
    new_n_n574_, new_n_n565_, new_n_n530_, new_n_n521_, new_n_n512_,
    new_n_n503_, new_n_n494_, new_n_n485_, new_n_n476_, new_n_n467_,
    new_n_n440_, new_n_n431_, new_n_n422_, new_n_n413_, new_n_n404_,
    new_n_n395_, new_n_n386_, new_n_n377_, new_n_n368_, new_n_n350_,
    new_n_n341_, new_n_n332_, new_n_n323_, new_n_n314_, new_n_n305_,
    new_n_n296_, new_n_n287_, new_n_n278_, new_n_n269_, new_n_n251_,
    new_n_n242_, new_n_n233_, new_n_n224_, new_n_n215_, new_n_n206_,
    new_n_n197_, new_n_n188_, new_n_n179_, new_n_n152_, new_n_n143_,
    new_n_n134_, new_n_n125_, new_n_n116_, new_n_n107_, new_n_n98_,
    new_n_n89_, new_n_n4_, new_n_n54_, new_n_n43_, new_ny0_, new_nj1_,
    new_nu1_, new_n_n55_, new_n_n42_, new_nx0_, new_nk1_, new_nt1_,
    new_n_n56_, new_n_n41_, new_na1_, new_nh1_, new_ns1_, new_n_n57_,
    new_n_n40_, new_nz0_, new_ni1_, new_nr1_, new_n_n0_, new_n_n877_,
    new_n_n866_, new_n_n768_, new_n_n58_, new_nb2_, new_n_n32_, new_n_n21_,
    new_n_n10_, new_n_n876_, new_n_n867_, new_n_n778_, new_n_n59_,
    new_nc2_, new_n_n33_, new_n_n20_, new_n_n11_, new_n_n897_, new_n_n886_,
    new_no0_, new_nd2_, new_n_n30_, new_n_n23_, new_n_n12_, new_n_n896_,
    new_n_n887_, new_n_n797_, new_ne2_, new_n_n31_, new_n_n22_, new_n_n13_,
    new_n_n1020_, new_n_n1009_, new_n_n998_, new_n_n917_, new_n_n906_,
    new_n_n807_, new_nb1_, new_nm1_, new_nx1_, new_ni2_, new_n_n25_,
    new_n_n14_, new_nn0_, new_n_n1021_, new_n_n1008_, new_n_n999_,
    new_n_n916_, new_n_n907_, new_n_n817_, new_nc1_, new_nl1_, new_ny1_,
    new_nh2_, new_n_n24_, new_n_n15_, new_n_n1029_, new_n_n1018_,
    new_n_n1011_, new_n_n1000_, new_n_n937_, new_n_n926_, new_n_n827_,
    new_n_n49_, new_n_n38_, new_nz1_, new_n_n34_, new_n_n27_, new_n_n16_,
    new_n_n1028_, new_n_n1019_, new_n_n1010_, new_n_n1001_, new_n_n936_,
    new_n_n927_, new_n_n837_, new_n_n48_, new_n_n39_, new_na2_, new_nj2_,
    new_n_n26_, new_n_n17_, new_n_n991_, new_n_n980_, new_n_n969_,
    new_n_n958_, new_n_n957_, new_n_n946_, new_n_n847_, new_n_n50_,
    new_n_n47_, new_n_n36_, new_nf1_, new_nq1_, new_n_n29_, new_n_n18_,
    new_n_n990_, new_n_n981_, new_n_n968_, new_n_n959_, new_n_n956_,
    new_n_n947_, new_n_n857_, new_n_n51_, new_n_n46_, new_n_n37_, new_ng1_,
    new_np1_, new_n_n28_, new_n_n19_, new_n_n989_, new_n_n978_,
    new_n_n971_, new_n_n960_, new_n_n52_, new_n_n45_, new_nw0_, new_nd1_,
    new_no1_, new_nv1_, new_ng2_, new_n_n988_, new_n_n979_, new_n_n970_,
    new_n_n961_, new_n_n53_, new_n_n44_, new_n_n35_, new_ne1_, new_nn1_,
    new_nw1_, new_nf2_;
  assign new_na0_ = pa0;
  assign new_nq_ = pq;
  assign new_nb0_ = pb0;
  assign new_nr_ = pr;
  assign new_nc0_ = pc0;
  assign new_ns_ = ps;
  assign new_nd0_ = pd0;
  assign new_nt_ = pt;
  assign new_ne0_ = pe0;
  assign new_nu_ = pu;
  assign new_nf0_ = pf0;
  assign new_nv_ = pv;
  assign new_ng0_ = pg0;
  assign new_nw_ = pw;
  assign new_nh0_ = ph0;
  assign new_nx_ = px;
  assign new_ni0_ = pi0;
  assign new_ny_ = py;
  assign new_nj0_ = pj0;
  assign new_nz_ = pz;
  assign new_nk0_ = pk0;
  assign new_nl0_ = pl0;
  assign new_nm0_ = pm0;
  assign pn0 = new_nn0_;
  assign po0 = new_no0_;
  assign pp0 = new_np0_;
  assign new_na_ = pa;
  assign new_nb_ = pb;
  assign new_nc_ = pc;
  assign new_nd_ = pd;
  assign new_ne_ = pe;
  assign new_nf_ = pf;
  assign new_ng_ = pg;
  assign new_nh_ = ph;
  assign new_ni_ = pi;
  assign new_nj_ = pj;
  assign new_nk_ = pk;
  assign new_nl_ = pl;
  assign new_nm_ = pm;
  assign new_nn_ = pn;
  assign new_no_ = po;
  assign new_n_n1017_ = new_no_ & new_n_n29_ & new_n_n26_ & new_n_n25_ & new_nh0_ & new_n_n27_ & new_n_n22_ & new_n_n20_ & new_n_n24_ & new_n_n30_;
  assign new_n_n1006_ = new_ni0_ & new_nd0_ & new_n_n30_ & new_n_n18_ & new_n_n21_ & new_nu_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n27_;
  assign new_n_n995_ = new_nv_ & new_nj0_ & new_n_n23_ & new_n_n21_ & new_nh0_ & new_nz_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n22_;
  assign new_n_n984_ = new_n_n27_ & new_n_n28_ & new_nj0_ & new_n_n22_ & new_nv_ & new_nf0_ & new_n_n21_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n32_ & new_n_n31_;
  assign new_n_n973_ = new_ni0_ & new_n_n27_ & new_n_n30_ & new_nv_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n28_;
  assign new_n_n962_ = new_nd_ & new_n_n27_ & new_n_n30_ & new_n_n5_ & new_n_n29_ & new_nf0_ & new_nk_ & new_n_n23_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n953_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_nk0_ & new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n32_;
  assign new_n_n942_ = new_n_n20_ & new_n_n27_ & new_nk0_ & new_ni0_ & new_n_n24_ & new_n_n23_ & new_n_n30_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n931_ = new_nk0_ & new_n_n27_ & new_n_n30_ & new_n_n18_ & new_n_n29_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n28_;
  assign new_n_n920_ = new_n_n27_ & new_n_n28_ & new_nd_ & new_ni0_ & new_n_n5_ & new_n_n30_ & new_nv_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n909_ = new_n_n28_ & new_n_n31_ & new_nk0_ & new_n_n27_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n21_ & new_n_n16_ & new_n_n10_ & new_n_n1_ & new_n_n33_ & new_n_n32_;
  assign new_n_n898_ = new_n_n15_ & new_n_n20_ & new_n_n30_ & new_nk0_ & new_n_n29_ & new_n_n25_ & new_n_n21_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n854_ = new_n_n28_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nk0_ & new_n_n25_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n34_ & new_n_n33_;
  assign new_n_n843_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nk0_ & new_ni0_ & new_n_n20_ & new_n_n21_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n832_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n15_ & new_ni0_ & new_n_n20_ & new_n_n2_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n821_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n29_ & new_n_n30_ & new_nk0_ & new_n_n15_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n810_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n28_ & new_n_n31_ & new_nj0_ & new_n_n22_ & new_n_n20_ & new_n_n27_ & new_n_n5_ & new_nd_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n799_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n3_ & new_n_n15_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n788_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n15_ & new_nd0_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_nk0_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n34_;
  assign new_n_n756_ = new_n_n20_ & new_n_n27_ & new_n_n21_ & new_nj0_ & new_n_n22_ & new_nf0_ & new_nh_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n745_ = new_n_n24_ & new_nl0_ & new_ni0_ & new_n_n21_ & new_n_n26_ & new_n_n25_ & new_n_n1_ & new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n20_;
  assign new_n_n734_ = new_n_n20_ & new_n_n27_ & new_ni0_ & new_nh0_ & new_n_n23_ & new_nz_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n28_;
  assign new_n_n723_ = new_n_n20_ & new_n_n27_ & new_n_n15_ & new_nl0_ & new_n_n21_ & new_n_n23_ & new_ni0_ & new_n_n26_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n28_;
  assign new_n_n712_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_n_n15_ & new_nl0_ & new_n_n26_ & new_n_n21_ & new_n_n0_ & new_n_n33_ & new_n_n10_ & new_n_n32_ & new_n_n17_;
  assign new_n_n701_ = new_n_n27_ & new_n_n28_ & new_n_n14_ & new_n_n20_ & new_nl0_ & new_ni0_ & new_n_n15_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n30_;
  assign new_n_n690_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nl0_ & new_n_n14_ & new_n_n26_ & new_n_n15_ & new_n_n24_ & new_n_n0_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n17_;
  assign new_n_n679_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nj0_ & new_nl0_ & new_n_n23_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n657_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_n_n15_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n646_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n21_ & new_n_n24_ & new_nl0_ & new_n_n2_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n635_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n16_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n7_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n624_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n21_ & new_n_n24_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n613_ = new_n_n33_ & new_n_n4_ & new_n_n3_ & new_n_n32_ & new_n_n31_ & new_n_n28_ & new_n_n30_ & new_n_n15_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n602_ = new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_n_n24_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n2_ & new_n_n21_ & new_n_n15_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n591_ = new_n_n33_ & new_n_n34_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n7_ & new_n_n15_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n580_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n15_ & new_n_n5_ & new_nd_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n569_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n3_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n16_ & new_nj0_ & new_nl0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n558_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n24_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n14_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n548_ = new_n_n30_ & new_nx_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n537_ = new_ni0_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_no_ & new_nh0_;
  assign new_n_n526_ = new_nq_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_nf0_ & new_ni0_;
  assign new_n_n515_ = new_nb0_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_ne0_ & new_ni0_;
  assign new_n_n504_ = new_nb0_ & new_n_n27_ & new_nf0_ & new_nj0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n493_ = new_ni0_ & new_no_ & new_nn_ & new_n_n30_ & new_nw_ & new_n_n27_ & new_nf0_;
  assign new_n_n482_ = new_nr_ & new_nm_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_ne0_ & new_ni0_;
  assign new_n_n471_ = new_nr_ & new_nm_ & new_n_n27_ & new_nf0_ & new_nj0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n460_ = new_n_n10_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_nj0_ & new_nm0_;
  assign new_n_n449_ = new_n_n25_ & new_nm0_ & new_n_n20_ & new_n_n14_ & new_ni0_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_n_n15_;
  assign new_n_n438_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n20_ & new_n_n2_ & new_nj_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n427_ = new_n_n15_ & new_n_n26_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_nm_ & new_n_n10_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n416_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n10_ & new_nm0_ & new_n_n20_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n405_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n20_ & new_nt_ & new_ni0_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n27_;
  assign new_n_n394_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n383_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n20_ & new_n_n10_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n29_;
  assign new_n_n372_ = new_n_n15_ & new_n_n26_ & new_n_n10_ & new_nm0_ & new_nt_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n8_ & new_n_n27_;
  assign new_n_n361_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_nm0_;
  assign new_n_n339_ = new_nm0_ & new_n_n27_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n328_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n317_ = new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n9_ & new_n_n14_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n306_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_nm_ & new_nt_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n295_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_nt_ & new_n_n10_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n284_ = new_n_n25_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n15_;
  assign new_n_n273_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n24_ & new_n_n14_ & new_n_n9_ & new_n_n1_ & new_nk_ & new_nm_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n262_ = new_n_n24_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n2_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n29_;
  assign new_n_n229_ = new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n218_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_nd_ & new_n_n20_ & new_n_n1_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n207_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_nd_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n27_ & new_nj0_;
  assign new_n_n196_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n10_ & new_n_n25_ & new_nk_ & new_nm_ & new_n_n9_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n185_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n20_ & new_n_n11_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n29_ & new_n_n27_;
  assign new_n_n174_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n29_;
  assign new_n_n163_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n23_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n119_ = new_n_n29_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n108_ = new_n_n27_ & new_n_n8_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n97_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n7_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n86_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n75_ = new_n_n29_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n64_ = new_n_n8_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n1016_ = new_no_ & new_n_n29_ & new_n_n26_ & new_n_n25_ & new_nh0_ & new_n_n27_ & new_n_n24_ & new_n_n22_ & new_nv_ & new_n_n30_;
  assign new_n_n1007_ = new_n_n22_ & new_nd0_ & new_n_n18_ & new_nj0_ & new_n_n21_ & new_nu_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n27_;
  assign new_n_n994_ = new_n_n30_ & new_nv_ & new_n_n23_ & new_n_n21_ & new_nh0_ & new_nz_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_ni0_;
  assign new_n_n985_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n20_ & new_nj0_ & new_nf0_ & new_n_n21_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n32_ & new_n_n31_;
  assign new_n_n972_ = new_n_n30_ & new_n_n27_ & new_n_n21_ & new_n_n29_ & new_nk_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n28_;
  assign new_n_n963_ = new_n_n28_ & new_n_n31_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_nf0_ & new_nk_ & new_n_n23_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_;
  assign new_n_n952_ = new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n20_ & new_n_n24_ & new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n943_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_nk0_ & new_n_n23_ & new_n_n30_ & new_n_n26_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n31_;
  assign new_n_n930_ = new_n_n24_ & new_nk0_ & new_n_n30_ & new_n_n18_ & new_n_n29_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n921_ = new_n_n31_ & new_n_n3_ & new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n30_ & new_nv_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n32_;
  assign new_n_n908_ = new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nk0_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n21_ & new_n_n16_ & new_n_n33_ & new_n_n1_ & new_n_n32_ & new_n_n31_;
  assign new_n_n899_ = new_ni0_ & new_n_n20_ & new_nk0_ & new_n_n15_ & new_n_n30_ & new_n_n25_ & new_n_n21_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n853_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n15_ & new_ni0_ & new_n_n25_ & new_n_n21_ & new_n_n30_ & new_nk0_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n844_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n15_ & new_ni0_ & new_n_n20_ & new_n_n21_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n831_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nk0_ & new_ni0_ & new_n_n20_ & new_n_n2_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n822_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n15_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n34_;
  assign new_n_n809_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n3_ & new_n_n22_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nk0_ & new_nj0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n800_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_nd_ & new_nk0_ & new_n_n15_ & new_ni0_ & new_n_n30_ & new_n_n24_ & new_n_n5_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n779_ = new_nj0_ & new_n_n24_ & new_n_n26_ & new_n_n22_ & new_n_n25_ & new_n_n1_ & new_n_n20_ & new_n_n27_ & new_n_n14_ & new_nl0_;
  assign new_n_n755_ = new_n_n28_ & new_n_n30_ & new_ni0_ & new_n_n27_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_nu_ & new_n_n31_;
  assign new_n_n746_ = new_n_n24_ & new_nl0_ & new_ni0_ & new_n_n15_ & new_n_n26_ & new_n_n25_ & new_n_n31_ & new_n_n27_ & new_n_n30_ & new_n_n20_ & new_n_n14_;
  assign new_n_n733_ = new_nh0_ & new_n_n27_ & new_ni0_ & new_n_n21_ & new_n_n23_ & new_nz_ & new_n_n33_ & new_n_n31_ & new_nu_ & new_n_n30_ & new_n_n28_;
  assign new_n_n724_ = new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n20_ & new_n_n21_ & new_n_n23_ & new_ni0_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n30_;
  assign new_n_n711_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n15_ & new_n_n24_ & new_n_n26_ & new_n_n21_ & new_n_n0_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n31_;
  assign new_n_n702_ = new_n_n28_ & new_n_n30_ & new_n_n20_ & new_n_n27_ & new_n_n14_ & new_ni0_ & new_nl0_ & new_n_n26_ & new_n_n23_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n31_;
  assign new_n_n689_ = new_n_n31_ & new_n_n17_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n14_ & new_n_n27_ & new_n_n26_ & new_n_n23_ & new_nl0_ & new_n_n0_ & new_n_n10_ & new_n_n1_ & new_n_n34_ & new_n_n33_;
  assign new_n_n680_ = new_n_n28_ & new_n_n30_ & new_n_n20_ & new_n_n27_ & new_nl0_ & new_n_n15_ & new_n_n24_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n33_ & new_n_n31_;
  assign new_n_n656_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n20_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_nn_;
  assign new_n_n647_ = new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n16_ & new_n_n21_ & new_nl0_ & new_n_n20_ & new_n_n2_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n634_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_n_n7_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n34_;
  assign new_n_n625_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n31_ & new_n_n17_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n21_ & new_nl0_ & new_nd0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n612_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n15_ & new_n_n5_ & new_nd_ & new_nl0_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n603_ = new_n_n33_ & new_n_n6_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n2_ & new_n_n21_ & new_n_n15_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n590_ = new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n7_ & new_n_n15_ & new_n_n24_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n34_;
  assign new_n_n581_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n30_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n16_ & new_n_n15_ & new_nl0_ & new_n_n14_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n559_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n17_ & new_n_n24_ & new_n_n3_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n31_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n557_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n17_ & new_n_n15_ & new_n_n3_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n31_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n549_ = new_nw_ & new_n_n27_ & new_n_n30_ & new_nx_ & new_ni0_;
  assign new_n_n536_ = new_n_n22_ & new_nw_ & new_ne0_ & new_n_n27_ & new_nj0_ & new_nx_;
  assign new_n_n527_ = new_nq_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_ng0_ & new_ni0_;
  assign new_n_n514_ = new_nb0_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_ng0_ & new_ni0_;
  assign new_n_n505_ = new_nb0_ & new_n_n27_ & new_nj0_ & new_ng0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n492_ = new_ni0_ & new_n_n20_ & new_nn_ & new_n_n27_ & new_n_n30_ & new_ne0_ & new_no_;
  assign new_n_n483_ = new_nr_ & new_nm_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nd0_;
  assign new_n_n470_ = new_nm0_ & new_n_n24_ & new_n_n20_ & new_n_n1_ & new_n_n30_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n26_;
  assign new_n_n461_ = new_n_n1_ & new_n_n14_ & new_n_n22_ & new_n_n20_ & new_n_n27_ & new_n_n24_ & new_n_n26_ & new_nj0_ & new_nm0_;
  assign new_n_n459_ = new_n_n10_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n26_ & new_nm0_ & new_n_n14_;
  assign new_n_n437_ = new_n_n15_ & new_n_n24_ & new_n_n14_ & new_nm0_ & new_n_n20_ & new_n_n2_ & new_nj_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n26_;
  assign new_n_n428_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_nm_ & new_n_n10_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n415_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n10_ & new_n_n14_ & new_n_n20_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n406_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n20_ & new_nt_ & new_ni0_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n393_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_nm0_;
  assign new_n_n384_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n20_ & new_n_n10_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n8_;
  assign new_n_n371_ = new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n14_ & new_nt_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n27_ & new_n_n26_;
  assign new_n_n362_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n338_ = new_n_n24_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n329_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n11_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n316_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n9_ & new_n_n10_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n307_ = new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_nm_ & new_n_n10_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n19_;
  assign new_n_n294_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n11_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n285_ = new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_n_n15_;
  assign new_n_n272_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n26_ & new_n_n1_ & new_n_n9_ & new_n_n10_ & new_nk_ & new_nm_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n263_ = new_nm0_ & new_n_n27_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n2_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n239_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n217_ = new_n_n24_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_nd_ & new_n_n20_ & new_n_n1_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n208_ = new_nm0_ & new_nj0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_nd_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n195_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n10_ & new_n_n14_ & new_nk_ & new_nm_ & new_n_n9_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n186_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n20_ & new_n_n11_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n29_;
  assign new_n_n173_ = new_n_n15_ & new_n_n24_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n29_ & new_n_n27_;
  assign new_n_n164_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n23_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n118_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n109_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n96_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n87_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n74_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n65_ = new_n_n27_ & new_n_n30_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n1026_ = new_n_n26_ & new_n_n25_ & new_nz_ & new_nh0_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_n_n24_ & new_nv_;
  assign new_n_n993_ = new_nd0_ & new_n_n27_ & new_n_n30_ & new_n_n18_ & new_n_n29_ & new_na_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n982_ = new_n_n27_ & new_n_n28_ & new_nv_ & new_ni0_ & new_n_n30_ & new_nf0_ & new_n_n21_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n32_ & new_n_n31_;
  assign new_n_n975_ = new_n_n22_ & new_n_n27_ & new_nv_ & new_nj0_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n28_;
  assign new_n_n964_ = new_n_n27_ & new_n_n28_ & new_nv_ & new_ni0_ & new_n_n30_ & new_nk_ & new_n_n21_ & new_nf0_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n31_;
  assign new_n_n955_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n30_ & new_nk0_ & new_n_n26_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n32_;
  assign new_n_n944_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_nk0_ & new_n_n23_ & new_n_n24_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n929_ = new_n_n3_ & new_n_n32_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n18_ & new_nd0_ & new_n_n29_ & new_n_n30_ & new_nc_ & new_n_n4_ & new_n_n6_ & new_n_n34_ & new_n_n33_;
  assign new_n_n918_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_nd_ & new_nk_ & new_n_n5_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n911_ = new_n_n31_ & new_n_n32_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n30_ & new_n_n18_ & new_n_n26_ & new_n_n29_ & new_n_n16_ & new_n_n10_ & new_n_n1_ & new_n_n34_ & new_n_n33_;
  assign new_n_n900_ = new_nk0_ & new_n_n15_ & new_n_n18_ & new_n_n24_ & new_n_n30_ & new_n_n25_ & new_n_n29_ & new_n_n26_ & new_n_n23_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n856_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nk0_ & new_n_n15_ & new_n_n25_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n34_;
  assign new_n_n845_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n28_ & new_n_n31_ & new_nk0_ & new_ni0_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n830_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n24_ & new_nk0_ & new_n_n15_ & new_ni0_ & new_n_n2_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n819_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n15_ & new_n_n27_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_nk0_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n812_ = new_n_n31_ & new_n_n32_ & new_n_n27_ & new_n_n28_ & new_n_n15_ & new_n_n24_ & new_nk0_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n33_;
  assign new_n_n801_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nd_ & new_nk0_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n24_ & new_n_n5_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n769_ = new_nd0_ & new_n_n27_ & new_n_n23_ & new_ni0_ & new_nv_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n28_;
  assign new_n_n758_ = new_n_n27_ & new_n_n28_ & new_nj0_ & new_n_n20_ & new_n_n22_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n747_ = new_nl0_ & new_n_n14_ & new_ni0_ & new_n_n24_ & new_n_n26_ & new_n_n25_ & new_n_n1_ & new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n20_;
  assign new_n_n732_ = new_nh0_ & new_n_n27_ & new_n_n22_ & new_nj0_ & new_n_n23_ & new_nz_ & new_n_n34_ & new_nu_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n721_ = new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n20_ & new_n_n24_ & new_n_n26_ & new_n_n21_ & new_nf0_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n29_;
  assign new_n_n714_ = new_n_n31_ & new_n_n17_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nl0_ & new_n_n27_ & new_n_n26_ & new_n_n21_ & new_n_n0_ & new_n_n10_ & new_n_n1_ & new_n_n33_ & new_n_n32_;
  assign new_n_n703_ = new_n_n28_ & new_n_n29_ & new_nl0_ & new_n_n27_ & new_n_n24_ & new_n_n21_ & new_n_n15_ & new_n_n26_ & new_n_n23_ & new_n_n0_ & new_n_n17_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n670_ = new_n_n31_ & new_n_n32_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n24_ & new_nl0_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_nj0_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n33_;
  assign new_n_n659_ = new_n_n33_ & new_n_n34_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n14_ & new_n_n20_ & new_n_n22_ & new_n_n16_ & new_nj0_ & new_nl0_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n648_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n2_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n33_;
  assign new_n_n633_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n15_ & new_nl0_ & new_n_n14_ & new_n_n7_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n34_;
  assign new_n_n622_ = new_n_n33_ & new_nn_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n615_ = new_n_n33_ & new_n_n4_ & new_n_n3_ & new_n_n32_ & new_n_n31_ & new_n_n28_ & new_n_n30_ & new_n_n24_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n604_ = new_n_n33_ & new_n_n6_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n2_ & new_n_n21_ & new_n_n24_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n589_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_n_n4_ & new_n_n32_ & new_n_n17_ & new_n_n3_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n31_ & new_n_n21_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n571_ = new_n_n33_ & new_n_n34_ & new_n_n3_ & new_n_n32_ & new_n_n31_ & new_n_n28_ & new_n_n30_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n16_ & new_n_n15_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n4_;
  assign new_n_n560_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n5_ & new_n_n17_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_nd_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n535_ = new_n_n22_ & new_nw_ & new_ng0_ & new_n_n27_ & new_nj0_ & new_nx_;
  assign new_n_n524_ = new_nq_ & new_n_n30_ & new_ng0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n517_ = new_nq_ & new_n_n27_ & new_nf0_ & new_nj0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n506_ = new_nb0_ & new_n_n27_ & new_nj0_ & new_ne0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n491_ = new_ni0_ & new_n_n20_ & new_nn_ & new_n_n27_ & new_n_n30_ & new_ng0_ & new_no_;
  assign new_n_n480_ = new_nr_ & new_nm_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_nf0_ & new_ni0_;
  assign new_n_n473_ = new_nr_ & new_nm_ & new_n_n27_ & new_nj0_ & new_ne0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n462_ = new_n_n1_ & new_nm0_ & new_n_n22_ & new_n_n20_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nj0_;
  assign new_n_n436_ = new_n_n15_ & new_n_n26_ & new_n_n10_ & new_nm0_ & new_n_n20_ & new_n_n2_ & new_nj_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n425_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n2_ & new_n_n14_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n418_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n20_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n407_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n20_ & new_n_n10_ & new_ni0_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n392_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_ni0_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_nm0_;
  assign new_n_n381_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n29_ & new_n_n27_;
  assign new_n_n374_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_nt_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n8_ & new_n_n27_;
  assign new_n_n363_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nm0_;
  assign new_n_n337_ = new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n326_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n319_ = new_n_n14_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_n_n15_ & new_nm0_;
  assign new_n_n308_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_nm_ & new_n_n10_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n19_;
  assign new_n_n293_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n11_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n282_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_n_n1_ & new_nm0_ & new_nk_ & new_nm_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n275_ = new_n_n26_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n1_ & new_nt_ & new_n_n10_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n29_;
  assign new_n_n264_ = new_n_n27_ & new_n_n29_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n2_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n238_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n20_ & new_n_n3_ & new_n_n1_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n227_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n209_ = new_nm0_ & new_nj0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_nd_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n27_ & new_n_n24_;
  assign new_n_n194_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_nt_ & new_n_n25_ & new_nk_ & new_nm_ & new_n_n9_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n183_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n29_ & new_n_n27_;
  assign new_n_n176_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n7_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n165_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n23_ & new_n_n11_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n139_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n13_ & new_n_n14_ & new_nd_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n128_ = new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n95_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n84_ = new_n_n15_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n77_ = new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n66_ = new_n_n8_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n1027_ = new_n_n25_ & new_no_ & new_nh0_ & new_n_n26_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_n_n24_ & new_nv_;
  assign new_n_n992_ = new_n_n18_ & new_nd0_ & new_n_n29_ & new_n_n30_ & new_n_n21_ & new_na_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n27_;
  assign new_n_n983_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_nf0_ & new_n_n21_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n32_ & new_n_n31_;
  assign new_n_n974_ = new_n_n20_ & new_n_n27_ & new_n_n30_ & new_ni0_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n28_;
  assign new_n_n965_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_nk_ & new_n_n21_ & new_nf0_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n31_;
  assign new_n_n954_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_nk0_ & new_n_n30_ & new_n_n24_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n945_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n20_ & new_nj0_ & new_n_n23_ & new_nk0_ & new_n_n26_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n31_;
  assign new_n_n928_ = new_n_n28_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_nd_ & new_n_n18_ & new_n_n5_ & new_n_n29_ & new_n_n30_ & new_nc_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n919_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_n_n22_ & new_nk_ & new_nj0_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_;
  assign new_n_n910_ = new_n_n28_ & new_n_n31_ & new_nk0_ & new_n_n27_ & new_n_n24_ & new_n_n30_ & new_n_n18_ & new_n_n26_ & new_n_n29_ & new_n_n16_ & new_n_n34_ & new_n_n1_ & new_n_n33_ & new_n_n32_;
  assign new_n_n901_ = new_n_n15_ & new_n_n27_ & new_n_n18_ & new_nk0_ & new_n_n30_ & new_n_n25_ & new_n_n29_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n855_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_nk0_ & new_n_n15_ & new_n_n25_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n34_;
  assign new_n_n846_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n20_ & new_n_n21_ & new_n_n24_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n829_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_nk0_ & new_n_n15_ & new_n_n20_ & new_n_n2_ & new_n_n29_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n820_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n15_ & new_n_n20_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n34_;
  assign new_n_n811_ = new_n_n6_ & new_n_n10_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_ & new_n_n32_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n31_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n802_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n28_ & new_n_n31_ & new_n_n15_ & new_ni0_ & new_n_n20_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n759_ = new_n_n28_ & new_n_n31_ & new_nj0_ & new_n_n27_ & new_n_n22_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_nu_;
  assign new_n_n757_ = new_n_n27_ & new_n_n28_ & new_n_n21_ & new_nj0_ & new_n_n22_ & new_nf0_ & new_nh_ & new_n_n32_ & new_n_n33_ & new_nu_ & new_n_n31_;
  assign new_n_n748_ = new_nj0_ & new_n_n20_ & new_n_n22_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n731_ = new_nh0_ & new_n_n20_ & new_n_n22_ & new_nj0_ & new_n_n23_ & new_nz_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n722_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_nl0_ & new_n_n21_ & new_n_n23_ & new_n_n22_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n28_;
  assign new_n_n713_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_n_n24_ & new_nl0_ & new_n_n26_ & new_n_n21_ & new_n_n0_ & new_n_n33_ & new_n_n1_ & new_n_n32_ & new_n_n17_;
  assign new_n_n704_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n21_ & new_n_n15_ & new_n_n26_ & new_n_n23_ & new_n_n0_ & new_n_n33_ & new_n_n10_ & new_n_n17_ & new_n_n31_;
  assign new_n_n669_ = new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_n_n21_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n23_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n660_ = new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nl0_ & new_n_n14_ & new_ni0_ & new_n_n16_ & new_n_n15_ & new_n_n24_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n34_ & new_n_n33_;
  assign new_n_n658_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nl0_ & new_n_n14_ & new_n_n22_ & new_n_n16_ & new_nj0_ & new_n_n24_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n34_;
  assign new_n_n632_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_n_n14_ & new_n_n20_ & new_n_n16_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n7_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n34_ & new_n_n33_;
  assign new_n_n623_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n21_ & new_n_n15_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n614_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_nl0_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n605_ = new_n_n6_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n2_ & new_n_n21_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n579_ = new_n_n33_ & new_n_n34_ & new_n_n3_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n16_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n4_;
  assign new_n_n570_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n14_ & new_ni0_ & new_n_n16_ & new_n_n15_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n34_;
  assign new_n_n561_ = new_n_n6_ & new_n_n10_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_ & new_nl0_ & new_n_n32_ & new_n_n29_ & new_n_n30_ & new_n_n31_ & new_n_n17_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n534_ = new_n_n22_ & new_nw_ & new_nj0_ & new_n_n27_ & new_nx_ & new_nf0_;
  assign new_n_n525_ = new_nq_ & new_n_n30_ & new_ne0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n516_ = new_nb0_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nd0_;
  assign new_n_n507_ = new_nb0_ & new_nw_ & new_nj0_ & new_n_n27_ & new_nf0_ & new_n_n22_;
  assign new_n_n490_ = new_ni0_ & new_n_n20_ & new_nn_ & new_n_n27_ & new_n_n30_ & new_nf0_ & new_no_;
  assign new_n_n481_ = new_nr_ & new_nm_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_ng0_ & new_ni0_;
  assign new_n_n472_ = new_nr_ & new_nm_ & new_n_n27_ & new_nj0_ & new_ng0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n463_ = new_n_n10_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n14_;
  assign new_n_n435_ = new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n14_ & new_n_n20_ & new_n_n2_ & new_nj_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n26_;
  assign new_n_n426_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n2_ & new_nm0_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n417_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n20_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n408_ = new_n_n27_ & new_n_n8_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n20_ & new_n_n10_ & new_ni0_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n391_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_ni0_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_nm0_ & new_n_n14_;
  assign new_n_n382_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n8_ & new_n_n29_;
  assign new_n_n373_ = new_n_n15_ & new_n_n24_ & new_n_n14_ & new_nm0_ & new_nt_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n27_ & new_n_n26_;
  assign new_n_n364_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n336_ = new_nm0_ & new_n_n27_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n327_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n318_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_n_n15_ & new_n_n24_ & new_n_n9_ & new_nm0_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n309_ = new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_nm_ & new_n_n14_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n19_;
  assign new_n_n292_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n283_ = new_n_n14_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_n_n15_ & new_nm0_;
  assign new_n_n274_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n9_ & new_n_n1_ & new_nk_ & new_nm_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n265_ = new_n_n24_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n1_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n237_ = new_n_n24_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n20_ & new_n_n3_ & new_n_n1_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n228_ = new_nm0_ & new_n_n27_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n219_ = new_n_n27_ & new_n_n29_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_nd_ & new_n_n10_ & new_n_n1_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n193_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_nt_ & new_n_n14_ & new_nk_ & new_nm_ & new_n_n9_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n184_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n29_;
  assign new_n_n175_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n7_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n166_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n23_ & new_n_n11_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n138_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n25_ & new_nd_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n129_ = new_n_n30_ & new_n_n19_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n14_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n94_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n85_ = new_n_n15_ & new_n_n24_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n27_;
  assign new_n_n76_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n67_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n1024_ = new_n_n24_ & new_nk0_ & new_n_n25_ & new_n_n30_ & new_n_n26_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n15_;
  assign new_n_n1013_ = new_n_n28_ & new_n_n31_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n1002_ = new_n_n18_ & new_ni0_ & new_n_n21_ & new_n_n30_ & new_n_n23_ & new_nu_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nd0_;
  assign new_n_n977_ = new_n_n27_ & new_n_n28_ & new_nv_ & new_ni0_ & new_n_n30_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n31_;
  assign new_n_n966_ = new_n_n27_ & new_n_n28_ & new_nj0_ & new_n_n22_ & new_nv_ & new_nk_ & new_n_n21_ & new_nf0_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n31_;
  assign new_n_n949_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_nk0_ & new_n_n21_ & new_n_n30_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n32_ & new_n_n31_;
  assign new_n_n938_ = new_nk0_ & new_n_n27_ & new_n_n18_ & new_n_n24_ & new_n_n30_ & new_n_n23_ & new_n_n29_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n935_ = new_n_n20_ & new_n_n27_ & new_nk0_ & new_ni0_ & new_n_n30_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n28_;
  assign new_n_n924_ = new_n_n27_ & new_n_n28_ & new_nj0_ & new_n_n22_ & new_nd_ & new_nv_ & new_n_n5_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n913_ = new_n_n28_ & new_n_n31_ & new_ni0_ & new_n_n27_ & new_nv_ & new_nk_ & new_n_n30_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_;
  assign new_n_n902_ = new_n_n20_ & new_n_n27_ & new_nk0_ & new_n_n15_ & new_n_n30_ & new_n_n25_ & new_n_n29_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n850_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nk0_ & new_n_n25_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n33_;
  assign new_n_n839_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_n_n18_ & new_nk0_ & new_nd0_ & new_n_n21_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n836_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n15_ & new_nd0_ & new_n_n30_ & new_n_n18_ & new_n_n24_ & new_nk0_ & new_n_n21_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_nn_;
  assign new_n_n825_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n30_ & new_n_n18_ & new_n_n24_ & new_nk0_ & new_n_n2_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n814_ = new_n_n31_ & new_n_n32_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nk0_ & new_n_n15_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n33_;
  assign new_n_n803_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n3_ & new_ni0_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n752_ = new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n28_;
  assign new_n_n741_ = new_n_n28_ & new_n_n30_ & new_nh0_ & new_n_n27_ & new_ni0_ & new_nz_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_nu_ & new_n_n31_;
  assign new_n_n738_ = new_n_n27_ & new_n_n28_ & new_nj0_ & new_nh0_ & new_n_n22_ & new_nz_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_nu_ & new_n_n31_;
  assign new_n_n727_ = new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n20_ & new_n_n15_ & new_ni0_ & new_n_n21_ & new_n_n26_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n716_ = new_n_n24_ & new_nl0_ & new_n_n21_ & new_nj0_ & new_n_n22_ & new_n_n26_ & new_n_n23_ & new_nf0_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n20_;
  assign new_n_n705_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n21_ & new_n_n24_ & new_n_n26_ & new_n_n23_ & new_n_n0_ & new_n_n33_ & new_n_n1_ & new_n_n17_ & new_n_n31_;
  assign new_n_n653_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n15_ & new_nl0_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n642_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_n_n16_ & new_n_n21_ & new_nj0_ & new_n_n24_ & new_n_n2_ & new_n_n22_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n628_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n23_ & new_n_n24_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n617_ = new_n_n4_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n30_ & new_n_n31_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n606_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_nj0_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n554_ = new_n_n33_ & new_n_n34_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n15_ & new_n_n30_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n544_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ne0_ & new_nb0_;
  assign new_n_n519_ = new_nq_ & new_n_n27_ & new_nj0_ & new_ne0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n508_ = new_nb0_ & new_nw_ & new_ng0_ & new_n_n27_ & new_nj0_ & new_n_n22_;
  assign new_n_n456_ = new_n_n26_ & new_n_n27_ & new_n_n1_ & new_nm0_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n445_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n14_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n409_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n20_ & new_n_n14_ & new_ni0_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n390_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n27_ & new_n_n8_ & new_n_n24_ & new_nj0_;
  assign new_n_n357_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n24_ & new_n_n27_ & new_nj0_ & new_nm0_;
  assign new_n_n346_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_n_n15_ & new_n_n24_ & new_nt_ & new_nm0_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n291_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n280_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n10_ & new_n_n1_ & new_nk_ & new_nm_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n258_ = new_nm0_ & new_n_n24_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n247_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n13_ & new_n_n14_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n192_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_nt_ & new_n_n10_ & new_nk_ & new_nm_ & new_n_n9_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n181_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n27_ & new_n_n24_;
  assign new_n_n170_ = new_n_n15_ & new_n_n24_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n2_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n27_;
  assign new_n_n159_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n2_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n29_ & new_n_n27_;
  assign new_n_n148_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_n_n3_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n93_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n82_ = new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_nm0_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n71_ = new_n_n29_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n60_ = new_n_n27_ & new_n_n8_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n9_ = ~new_nd_;
  assign new_n_n1025_ = new_n_n24_ & new_nk0_ & new_n_n25_ & new_n_n30_ & new_n_n26_ & new_n_n1_ & new_n_n27_ & new_n_n31_ & new_n_n20_ & new_ni0_;
  assign new_n_n1012_ = new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n21_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n32_ & new_n_n31_;
  assign new_n_n1003_ = new_nj0_ & new_n_n22_ & new_n_n21_ & new_n_n18_ & new_n_n23_ & new_nu_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nd0_;
  assign new_n_n976_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n28_;
  assign new_n_n967_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n20_ & new_nj0_ & new_nk_ & new_n_n21_ & new_nf0_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n31_;
  assign new_n_n948_ = new_n_n20_ & new_n_n27_ & new_nk0_ & new_ni0_ & new_n_n24_ & new_n_n21_ & new_n_n30_ & new_n_n26_ & new_n_n1_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n939_ = new_n_n27_ & new_n_n28_ & new_n_n18_ & new_nk0_ & new_n_n30_ & new_n_n23_ & new_n_n29_ & new_n_n26_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n31_;
  assign new_n_n934_ = new_ni0_ & new_n_n20_ & new_n_n24_ & new_nk0_ & new_n_n30_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n925_ = new_n_n31_ & new_n_n3_ & new_n_n27_ & new_n_n28_ & new_n_n22_ & new_nv_ & new_nj0_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n32_;
  assign new_n_n912_ = new_ni0_ & new_n_n27_ & new_n_n5_ & new_nd_ & new_nv_ & new_nk_ & new_n_n30_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n903_ = new_n_n20_ & new_n_n27_ & new_n_n15_ & new_ni0_ & new_nk0_ & new_n_n25_ & new_n_n30_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n849_ = new_n_n28_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n15_ & new_n_n18_ & new_nk0_ & new_n_n25_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n33_;
  assign new_n_n840_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n15_ & new_n_n21_ & new_n_n29_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n835_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n28_ & new_n_n31_ & new_nj0_ & new_n_n22_ & new_n_n20_ & new_n_n27_ & new_n_n2_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n826_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n30_ & new_n_n18_ & new_nk0_ & new_n_n15_ & new_n_n2_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n813_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nk0_ & new_n_n15_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n804_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n15_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n5_ & new_nd_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n751_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_nj0_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_nu_ & new_n_n31_;
  assign new_n_n742_ = new_n_n15_ & new_n_n24_ & new_n_n22_ & new_n_n21_ & new_n_n26_ & new_n_n25_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n20_ & new_nl0_;
  assign new_n_n737_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_nh0_ & new_n_n22_ & new_nz_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n728_ = new_n_n28_ & new_n_n30_ & new_n_n20_ & new_n_n27_ & new_nl0_ & new_ni0_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n32_ & new_n_n31_;
  assign new_n_n715_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nl0_ & new_n_n14_ & new_n_n26_ & new_n_n15_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n706_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_n_n21_ & new_nl0_ & new_n_n26_ & new_n_n23_ & new_n_n0_ & new_n_n10_ & new_n_n1_ & new_n_n33_ & new_n_n17_;
  assign new_n_n652_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_nn_;
  assign new_n_n643_ = new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n21_ & new_nj0_ & new_nl0_ & new_n_n2_ & new_n_n22_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n638_ = new_n_n17_ & new_n_n32_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_nd0_ & new_n_n7_ & new_n_n21_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n33_;
  assign new_n_n616_ = new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n607_ = new_n_n33_ & new_n_n4_ & new_n_n3_ & new_n_n32_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nj0_ & new_n_n24_ & new_nl0_ & new_n_n20_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_np0_ = new_n_n418_ | new_nn1_ | new_n_n400_ | new_n_n409_ | new_n_n382_ | new_n_n391_ | new_n_n348_ | new_n_n373_ | new_n_n330_ | new_n_n339_ | new_n_n312_ | new_n_n321_ | new_n_n294_ | new_n_n303_ | new_n_n276_ | new_n_n285_ | new_n_n251_ | new_n_n260_ | new_n_n233_ | new_n_n242_ | new_n_n215_ | new_n_n224_ | new_n_n197_ | new_n_n206_ | new_n_n154_ | new_n_n163_ | new_n_n136_ | new_n_n145_ | new_n_n66_ | new_n_n127_ | new_n_n57_ | new_n_n419_ | new_nf1_ | new_n_n401_ | new_n_n408_ | new_n_n383_ | new_n_n390_ | new_n_n358_ | new_n_n372_ | new_n_n329_ | new_n_n340_ | new_n_n311_ | new_n_n322_ | new_n_n293_ | new_n_n304_ | new_n_n275_ | new_n_n286_ | new_n_n250_ | new_n_n261_ | new_n_n232_ | new_n_n243_ | new_n_n214_ | new_n_n225_ | new_n_n196_ | new_n_n207_ | new_n_n153_ | new_n_n164_ | new_n_n135_ | new_n_n146_ | new_n_n67_ | new_n_n117_ | new_nr1_ | new_n_n56_ | new_n_n438_ | new_n_n402_ | new_n_n429_ | new_n_n380_ | new_n_n393_ | new_n_n341_ | new_n_n371_ | new_n_n319_ | new_n_n332_ | new_n_n305_ | new_n_n310_ | new_n_n283_ | new_n_n296_ | new_n_n258_ | new_n_n274_ | new_n_n244_ | new_n_n249_ | new_n_n222_ | new_n_n235_ | new_n_n186_ | new_n_n213_ | new_n_n161_ | new_n_n177_ | new_n_n147_ | new_n_n152_ | new_n_n116_ | new_n_n125_ | new_n_n55_ | new_n_n64_ | new_n_n439_ | new_no1_ | new_n_n403_ | new_n_n428_ | new_n_n392_ | new_n_n370_ | new_n_n381_ | new_n_n331_ | new_n_n342_ | new_n_n309_ | new_n_n320_ | new_n_n295_ | new_n_n306_ | new_n_n273_ | new_n_n284_ | new_n_n248_ | new_n_n259_ | new_n_n234_ | new_n_n245_ | new_n_n212_ | new_n_n223_ | new_n_n187_ | new_n_n162_ | new_n_n176_ | new_n_n137_ | new_n_n151_ | new_n_n115_ | new_n_n126_ | new_n_n54_ | new_n_n65_ | new_n_n431_ | new_n_n440_ | new_n_n413_ | new_n_n422_ | new_n_n369_ | new_n_n378_ | new_n_n334_ | new_n_n343_ | new_n_n325_ | new_n_n299_ | new_n_n316_ | new_n_n281_ | new_n_n290_ | new_n_n246_ | new_n_n272_ | new_n_n202_ | new_n_n237_ | new_n_n184_ | new_n_n193_ | new_n_n159_ | new_n_n175_ | new_n_n105_ | new_n_n150_ | new_n_n87_ | new_n_n96_ | new_n_n53_ | new_n_n62_ | new_n_n441_ | new_ns1_ | new_n_n423_ | new_n_n430_ | new_n_n379_ | new_n_n412_ | new_n_n344_ | new_n_n368_ | new_n_n326_ | new_n_n333_ | new_n_n300_ | new_n_n315_ | new_n_n282_ | new_n_n289_ | new_n_n271_ | new_n_n236_ | new_n_n247_ | new_n_n192_ | new_n_n203_ | new_n_n174_ | new_n_n185_ | new_n_n149_ | new_n_n160_ | new_n_n95_ | new_n_n106_ | new_n_n63_ | new_n_n77_ | new_n_n442_ | new_n_n52_ | new_n_n420_ | new_n_n433_ | new_n_n398_ | new_n_n411_ | new_n_n345_ | new_n_n389_ | new_n_n323_ | new_n_n336_ | new_n_n301_ | new_n_n314_ | new_n_n279_ | new_n_n292_ | new_n_n226_ | new_n_n270_ | new_n_n204_ | new_n_n217_ | new_n_n182_ | new_n_n195_ | new_n_n173_ | new_n_n107_ | new_n_n148_ | new_n_n76_ | new_n_n85_ | new_n_n51_ | new_n_n60_ | new_n_n432_ | new_n_n443_ | new_n_n410_ | new_n_n421_ | new_n_n388_ | new_n_n399_ | new_n_n335_ | new_n_n346_ | new_n_n313_ | new_n_n324_ | new_n_n291_ | new_n_n302_ | new_n_n269_ | new_n_n280_ | new_n_n216_ | new_n_n227_ | new_n_n194_ | new_n_n205_ | new_n_n172_ | new_n_n183_ | new_n_n97_ | new_n_n158_ | new_n_n75_ | new_n_n86_ | new_n_n50_ | new_n_n61_ | new_n_n508_ | new_n_n490_ | new_n_n499_ | new_n_n472_ | new_n_n481_ | new_n_n435_ | new_n_n444_ | new_n_n417_ | new_n_n426_ | new_n_n58_ | new_n_n347_ | new_n_n509_ | new_n_n49_ | new_n_n491_ | new_n_n498_ | new_n_n473_ | new_n_n480_ | new_n_n445_ | new_n_n427_ | new_n_n434_ | new_n_n337_ | new_n_n416_ | new_n_n48_ | new_n_n59_ | new_n_n501_ | new_n_n510_ | new_n_n479_ | new_n_n488_ | new_n_n446_ | new_n_n474_ | new_n_n424_ | new_n_n437_ | new_n_n327_ | new_n_n415_ | new_n_n511_ | new_n_n489_ | new_n_n500_ | new_n_n475_ | new_n_n478_ | new_n_n436_ | new_n_n447_ | new_n_n414_ | new_n_n425_ | new_nu1_ | new_n_n317_ | new_n_n512_ | new_n_n547_ | new_n_n494_ | new_n_n503_ | new_n_n468_ | new_n_n485_ | new_n_n395_ | new_n_n404_ | new_n_n377_ | new_n_n386_ | new_nt1_ | new_n_n307_ | new_n_n513_ | new_n_n546_ | new_n_n495_ | new_n_n502_ | new_n_n469_ | new_n_n484_ | new_n_n394_ | new_n_n405_ | new_n_n376_ | new_n_n387_ | new_n_n297_ | new_n_n527_ | new_n_n536_ | new_n_n505_ | new_n_n514_ | new_n_n483_ | new_n_n492_ | new_n_n406_ | new_n_n470_ | new_n_n384_ | new_n_n397_ | new_n_n287_ | new_n_n375_ | new_n_n526_ | new_n_n537_ | new_n_n504_ | new_n_n515_ | new_n_n482_ | new_n_n493_ | new_n_n407_ | new_n_n471_ | new_n_n385_ | new_n_n396_ | new_n_n277_ | new_n_n374_ | new_n_n543_ | new_n_n552_ | new_n_n525_ | new_n_n534_ | new_n_n507_ | new_n_n516_ | new_n_n542_ | new_n_n553_ | new_n_n535_ | new_n_n517_ | new_n_n524_ | new_nz1_ | new_n_n506_ | new_n_n532_ | new_n_n545_ | new_n_n496_ | new_n_n523_ | new_nv1_ | new_n_n487_ | new_n_n533_ | new_n_n544_ | new_n_n497_ | new_n_n522_ | new_n_n548_ | new_n_n486_ | new_n_n530_ | new_n_n539_ | new_n_n476_ | new_n_n521_ | new_n_n457_ | new_n_n466_ | new_n_n538_ | new_n_n549_ | new_n_n520_ | new_n_n531_ | new_n_n467_ | new_n_n477_ | new_n_n550_ | new_n_n456_ | new_n_n528_ | new_n_n541_ | new_n_n519_ | new_n_n455_ | new_n_n464_ | new_n_n38_ | new_n_n367_ | new_n_n540_ | new_n_n551_ | new_n_n518_ | new_n_n529_ | new_n_n454_ | new_n_n465_ | new_n_n39_ | new_n_n357_ | new_n_n453_ | new_n_n462_ | new_n_n356_ | new_n_n365_ | new_n_n268_ | new_n_n189_ | new_n_n198_ | new_n_n171_ | new_n_n180_ | new_n_n119_ | new_n_n128_ | new_n_n101_ | new_n_n110_ | new_n_n83_ | new_n_n92_ | new_n_n40_ | new_n_n74_ | new_n_n452_ | new_n_n463_ | new_n_n355_ | new_n_n366_ | new_n_n278_ | new_n_n188_ | new_n_n199_ | new_n_n170_ | new_n_n181_ | new_n_n120_ | new_n_n138_ | new_n_n102_ | new_n_n109_ | new_n_n84_ | new_n_n91_ | new_n_n41_ | new_n_n73_ | new_n_n460_ | new_na1_ | new_n_n363_ | new_n_n451_ | new_n_n288_ | new_n_n354_ | new_n_n257_ | new_n_n266_ | new_n_n191_ | new_n_n200_ | new_n_n169_ | new_n_n178_ | new_n_n130_ | new_n_n139_ | new_n_n103_ | new_n_n108_ | new_n_n81_ | new_n_n94_ | new_n_n42_ | new_n_n72_ | new_n_n461_ | new_n_n364_ | new_n_n450_ | new_n_n298_ | new_n_n353_ | new_n_n256_ | new_n_n267_ | new_n_n190_ | new_n_n201_ | new_n_n168_ | new_n_n179_ | new_n_n129_ | new_n_n140_ | new_n_n104_ | new_n_n118_ | new_n_n82_ | new_n_n93_ | new_n_n71_ | new_nc1_ | new_n_n43_ | new_n_n449_ | new_n_n458_ | new_n_n352_ | new_n_n361_ | new_n_n264_ | new_n_n308_ | new_n_n238_ | new_n_n255_ | new_n_n220_ | new_n_n229_ | new_n_n167_ | new_n_n211_ | new_n_n132_ | new_n_n141_ | new_n_n123_ | new_n_n88_ | new_n_n114_ | new_n_n70_ | new_n_n79_ | new_n_n35_ | new_n_n44_ | new_n_n459_ | new_nb1_ | new_n_n362_ | new_n_n448_ | new_n_n318_ | new_n_n351_ | new_n_n254_ | new_n_n265_ | new_n_n228_ | new_n_n239_ | new_n_n210_ | new_n_n221_ | new_n_n142_ | new_n_n157_ | new_n_n124_ | new_n_n131_ | new_n_n98_ | new_n_n113_ | new_n_n69_ | new_n_n80_ | new_ne1_ | new_n_n45_ | new_n_n350_ | new_n_n359_ | new_n_n262_ | new_n_n328_ | new_n_n253_ | new_n_n231_ | new_n_n240_ | new_n_n209_ | new_n_n218_ | new_n_n156_ | new_n_n165_ | new_n_n134_ | new_n_n143_ | new_n_n112_ | new_n_n121_ | new_n_n90_ | new_n_n99_ | new_n_n46_ | new_n_n68_ | new_nd1_ | new_n_n37_ | new_n_n360_ | new_n_n338_ | new_n_n349_ | new_n_n252_ | new_n_n263_ | new_n_n230_ | new_n_n241_ | new_n_n208_ | new_n_n219_ | new_n_n155_ | new_n_n166_ | new_n_n133_ | new_n_n144_ | new_n_n111_ | new_n_n122_ | new_n_n89_ | new_n_n100_ | new_n_n78_ | new_n_n36_ | new_n_n47_;
  assign new_n_n545_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_nf0_ & new_nq_;
  assign new_n_n518_ = new_nq_ & new_n_n27_ & new_nj0_ & new_ng0_ & new_n_n20_ & new_n_n22_;
  assign new_n_n509_ = new_nb0_ & new_nw_ & new_ne0_ & new_n_n27_ & new_nj0_ & new_n_n22_;
  assign new_n_n455_ = new_nm0_ & new_n_n26_ & new_n_n1_ & new_n_n14_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n446_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n25_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n419_ = new_n_n15_ & new_n_n26_ & new_n_n14_ & new_nm0_ & new_n_n10_ & new_n_n2_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n380_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n8_ & new_n_n29_;
  assign new_n_n356_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_n_n22_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n27_ & new_n_n8_ & new_nj0_ & new_nm0_;
  assign new_n_n347_ = new_n_n27_ & new_n_n29_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n1_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n290_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n281_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n1_ & new_n_n14_ & new_nk_ & new_nm_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n257_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n27_ & new_n_n24_;
  assign new_n_n248_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n25_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n191_ = new_n_n15_ & new_n_n26_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_nt_ & new_n_n10_ & new_nk_ & new_nm_ & new_n_n9_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n182_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n160_ = new_n_n15_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n2_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n29_;
  assign new_n_n158_ = new_n_n15_ & new_n_n24_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n2_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n27_;
  assign new_n_n149_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n13_ & new_n_n14_ & new_n_n20_ & new_n_n3_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n92_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n83_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n27_;
  assign new_n_n70_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n61_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n1022_ = new_n_n30_ & new_n_n18_ & new_n_n26_ & new_n_n25_ & new_nu_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_ni0_ & new_n_n24_;
  assign new_n_n1015_ = new_n_n25_ & new_n_n30_ & new_nh0_ & new_n_n26_ & new_nz_ & new_n_n31_ & new_ni0_ & new_n_n27_ & new_n_n24_ & new_nv_;
  assign new_n_n1004_ = new_ni0_ & new_nd0_ & new_n_n30_ & new_n_n18_ & new_n_n23_ & new_nu_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n997_ = new_nj0_ & new_n_n22_ & new_n_n21_ & new_nv_ & new_nh0_ & new_nz_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n27_;
  assign new_n_n986_ = new_n_n28_ & new_n_n31_ & new_ni0_ & new_n_n27_ & new_nv_ & new_nf0_ & new_n_n30_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n951_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n20_ & new_nj0_ & new_n_n21_ & new_nk0_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n32_ & new_n_n31_;
  assign new_n_n940_ = new_n_n20_ & new_n_n27_ & new_n_n24_ & new_nk0_ & new_n_n30_ & new_n_n23_ & new_n_n29_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n933_ = new_n_n20_ & new_n_n27_ & new_n_n30_ & new_nk0_ & new_n_n29_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n28_;
  assign new_n_n922_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_nd_ & new_n_n30_ & new_n_n5_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n915_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_nk_ & new_n_n30_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_;
  assign new_n_n904_ = new_n_n20_ & new_n_n27_ & new_nk0_ & new_n_n15_ & new_n_n30_ & new_n_n21_ & new_n_n29_ & new_n_n26_ & new_n_n25_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n852_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_nk0_ & new_n_n15_ & new_n_n25_ & new_n_n21_ & new_n_n30_ & new_n_n24_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n33_;
  assign new_n_n841_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_nk0_ & new_n_n15_ & new_n_n20_ & new_n_n21_ & new_n_n29_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n834_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n20_ & new_n_n2_ & new_n_n24_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n823_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n30_ & new_nk0_ & new_n_n15_ & new_ni0_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n816_ = new_n_n31_ & new_n_n32_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n15_ & new_ni0_ & new_n_n21_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n33_;
  assign new_n_n805_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n28_ & new_n_n31_ & new_nk0_ & new_ni0_ & new_n_n20_ & new_n_n27_ & new_n_n30_ & new_n_n5_ & new_nd_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n754_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n30_;
  assign new_n_n743_ = new_n_n24_ & new_nl0_ & new_n_n22_ & new_n_n15_ & new_n_n26_ & new_n_n25_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n20_ & new_n_n14_;
  assign new_n_n736_ = new_nh0_ & new_n_n27_ & new_n_n21_ & new_nj0_ & new_n_n22_ & new_nz_ & new_n_n33_ & new_nu_ & new_n_n32_ & new_n_n31_ & new_n_n28_;
  assign new_n_n725_ = new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n20_ & new_n_n15_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n29_;
  assign new_n_n718_ = new_n_n20_ & new_n_n27_ & new_n_n24_ & new_nl0_ & new_n_n21_ & new_n_n26_ & new_n_n23_ & new_nf0_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n28_;
  assign new_n_n707_ = new_n_n28_ & new_n_n29_ & new_n_n20_ & new_n_n27_ & new_n_n14_ & new_n_n15_ & new_nl0_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n30_;
  assign new_n_n655_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_ & new_n_n30_ & new_n_n21_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n644_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_n_n2_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n33_;
  assign new_n_n637_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n15_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n34_;
  assign new_n_n626_ = new_n_n17_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n23_ & new_n_n15_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n34_;
  assign new_n_n608_ = new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n556_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n15_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n14_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n546_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ng0_ & new_nq_;
  assign new_n_n539_ = new_no_ & new_nn_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nf0_;
  assign new_n_n528_ = new_nq_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_ne0_ & new_ni0_;
  assign new_n_n458_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n24_ & new_n_n1_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n447_ = new_n_n14_ & new_n_n25_ & new_n_n20_ & new_n_n10_ & new_ni0_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_nm0_;
  assign new_n_n429_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_nm_ & new_n_n14_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n370_ = new_n_n24_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n359_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_ni0_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_nm0_ & new_n_n14_;
  assign new_n_n348_ = new_n_n29_ & new_n_n8_ & new_nm0_ & new_n_n27_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n1_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n271_ = new_n_n26_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n1_ & new_n_n9_ & new_n_n10_ & new_nk_ & new_nm_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n260_ = new_nm0_ & new_n_n27_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n2_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n29_;
  assign new_n_n249_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n14_ & new_n_n25_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n190_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n25_ & new_n_n2_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n172_ = new_n_n15_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n2_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n29_;
  assign new_n_n161_ = new_n_n15_ & new_n_n24_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n29_ & new_n_n27_;
  assign new_n_n91_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n80_ = new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n73_ = new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n62_ = new_n_n27_ & new_n_n8_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n1023_ = new_n_n30_ & new_n_n24_ & new_n_n25_ & new_n_n29_ & new_n_n26_ & new_n_n27_ & new_n_n22_ & new_n_n20_ & new_n_n15_ & new_nk0_;
  assign new_n_n1014_ = new_n_n25_ & new_n_n29_ & new_nh0_ & new_n_n26_ & new_nz_ & new_n_n27_ & new_n_n24_ & new_n_n22_ & new_nv_ & new_n_n30_;
  assign new_n_n1005_ = new_n_n22_ & new_nd0_ & new_n_n18_ & new_nj0_ & new_n_n23_ & new_nu_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n996_ = new_nv_ & new_ni0_ & new_n_n21_ & new_n_n30_ & new_nh0_ & new_nz_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n27_;
  assign new_n_n987_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_nf0_ & new_n_n30_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n950_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_nk0_ & new_n_n21_ & new_n_n24_ & new_n_n26_ & new_n_n1_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n941_ = new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n20_ & new_n_n30_ & new_n_n23_ & new_n_n29_ & new_n_n26_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n31_;
  assign new_n_n932_ = new_nk0_ & new_n_n20_ & new_n_n30_ & new_n_n24_ & new_n_n29_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n923_ = new_n_n31_ & new_n_n3_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n30_ & new_ni0_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n32_;
  assign new_n_n914_ = new_n_n20_ & new_n_n27_ & new_nd_ & new_ni0_ & new_n_n5_ & new_nk_ & new_n_n30_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n905_ = new_n_n20_ & new_n_n27_ & new_n_n15_ & new_ni0_ & new_nk0_ & new_n_n21_ & new_n_n30_ & new_n_n26_ & new_n_n25_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n851_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nk0_ & new_n_n15_ & new_n_n25_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n842_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n24_ & new_nk0_ & new_n_n15_ & new_ni0_ & new_n_n21_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n833_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n28_ & new_n_n31_ & new_nk0_ & new_ni0_ & new_n_n20_ & new_n_n27_ & new_n_n2_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n824_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n15_ & new_nd0_ & new_n_n30_ & new_n_n18_ & new_n_n24_ & new_nk0_ & new_n_n2_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n34_;
  assign new_n_n815_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n15_ & new_n_n20_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_nk0_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n806_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n3_ & new_ni0_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_nk0_ & new_n_n15_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n753_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_nu_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n744_ = new_n_n15_ & new_n_n24_ & new_ni0_ & new_n_n21_ & new_n_n26_ & new_n_n25_ & new_n_n31_ & new_n_n27_ & new_n_n30_ & new_n_n20_ & new_nl0_;
  assign new_n_n735_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_nh0_ & new_n_n23_ & new_nz_ & new_n_n34_ & new_nu_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n726_ = new_n_n27_ & new_n_n28_ & new_nl0_ & new_n_n20_ & new_nj0_ & new_n_n22_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n32_ & new_n_n31_;
  assign new_n_n717_ = new_nl0_ & new_n_n20_ & new_n_n21_ & new_n_n24_ & new_ni0_ & new_n_n26_ & new_n_n23_ & new_nf0_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n27_;
  assign new_n_n708_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_n_n14_ & new_nj0_ & new_nl0_ & new_n_n26_ & new_n_n22_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n32_;
  assign new_n_n654_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n24_ & new_nl0_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n645_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_nl0_ & new_n_n2_ & new_ni0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n636_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_n_n7_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n34_ & new_n_n33_;
  assign new_n_n627_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n23_ & new_n_n15_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n618_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n33_;
  assign new_n_n555_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n31_ & new_n_n15_ & new_n_n17_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n547_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ne0_ & new_nq_;
  assign new_n_n538_ = new_nd0_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nx_;
  assign new_n_n529_ = new_nq_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nd0_;
  assign new_n_n457_ = new_n_n24_ & new_n_n26_ & new_n_n14_ & new_nm0_ & new_n_n1_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n448_ = new_n_n25_ & new_nm0_ & new_n_n20_ & new_n_n10_ & new_ni0_ & new_n_n30_ & new_n_n27_ & new_n_n8_ & new_n_n26_ & new_n_n15_;
  assign new_n_n439_ = new_nm0_ & new_n_n26_ & new_n_n1_ & new_n_n14_ & new_n_n10_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n360_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_ni0_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_nm0_;
  assign new_n_n358_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n27_ & new_n_n8_ & new_n_n24_ & new_nj0_;
  assign new_n_n349_ = new_n_n30_ & new_n_n19_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n14_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n270_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n24_ & new_n_n1_ & new_n_n9_ & new_nt_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n261_ = new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n2_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n29_ & new_n_n27_;
  assign new_n_n259_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n2_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n29_ & new_n_n27_;
  assign new_n_n180_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n25_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n2_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n171_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n2_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n29_ & new_n_n27_;
  assign new_n_n162_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n29_;
  assign new_n_n90_ = new_n_n27_ & new_n_n8_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n81_ = new_n_n30_ & new_n_n19_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n14_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n72_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n63_ = new_n_n27_ & new_n_n30_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n895_ = new_n_n28_ & new_n_n31_ & new_n_n15_ & new_n_n27_ & new_nk0_ & new_n_n30_ & new_n_n18_ & new_n_n26_ & new_n_n25_ & new_n_n29_ & new_n_n16_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n32_;
  assign new_n_n884_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_n_n24_ & new_nk0_ & new_n_n23_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n34_;
  assign new_n_n873_ = new_n_n34_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_nk0_ & new_ni0_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n862_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nk0_ & new_n_n20_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n796_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n5_ & new_nd_ & new_nk0_ & new_n_n15_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n786_ = new_n_n26_ & new_n_n22_ & new_nz_ & new_n_n25_ & new_nu_ & new_nh0_ & new_n_n27_ & new_n_n24_ & new_nj0_;
  assign new_n_n775_ = new_ni0_ & new_n_n24_ & new_n_n25_ & new_n_n26_ & new_nz_ & new_nu_ & new_n_n30_ & new_n_n31_ & new_n_n27_ & new_nh0_;
  assign new_n_n764_ = new_n_n28_ & new_n_n29_ & new_nd0_ & new_n_n27_ & new_n_n21_ & new_nc_ & new_n_n33_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n30_;
  assign new_n_n698_ = new_n_n27_ & new_n_n28_ & new_n_n14_ & new_n_n20_ & new_nl0_ & new_ni0_ & new_n_n24_ & new_nf0_ & new_n_n26_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n687_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nl0_ & new_n_n14_ & new_n_n26_ & new_n_n23_ & new_n_n15_ & new_n_n0_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n17_;
  assign new_n_n676_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n33_ & new_n_n32_;
  assign new_n_n665_ = new_n_n31_ & new_n_n33_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n15_ & new_nl0_ & new_n_n14_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n34_;
  assign new_n_n649_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n15_ & new_nl0_ & new_n_n20_ & new_n_n2_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n588_ = new_n_n6_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n21_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n577_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n3_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_ni0_ & new_n_n16_ & new_nl0_ & new_n_n14_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n566_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n14_ & new_n_n22_ & new_n_n16_ & new_nj0_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n551_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_nx_ & new_nf0_;
  assign new_n_n540_ = new_no_ & new_nn_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_ng0_;
  assign new_n_n479_ = new_nr_ & new_nm_ & new_n_n30_ & new_ne0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n468_ = new_n_n1_ & new_nm0_ & new_n_n20_ & new_n_n10_ & new_n_n30_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n26_;
  assign new_n_n452_ = new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n25_ & new_n_n20_ & new_n_n30_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n26_;
  assign new_n_n441_ = new_n_n24_ & new_n_n26_ & new_n_n14_ & new_nm0_ & new_n_n1_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n430_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_nm_ & new_n_n25_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n369_ = new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n353_ = new_n_n30_ & new_n_n19_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_n_n15_ & new_n_n24_ & new_n_n14_ & new_nm0_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n342_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n20_ & new_n_n1_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n331_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n27_ & new_nj0_;
  assign new_n_n320_ = new_n_n25_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n15_;
  assign new_n_n254_ = new_nm0_ & new_nj0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n2_ & new_n_n22_ & new_n_n16_ & new_n_n8_ & new_n_n6_ & new_n_n27_ & new_n_n24_;
  assign new_n_n243_ = new_n_n27_ & new_n_n29_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n3_ & new_n_n10_ & new_n_n1_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n232_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n221_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n24_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_nd_ & new_n_n1_ & new_n_n11_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n210_ = new_nj0_ & new_n_n24_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_nd_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n155_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n27_ & new_n_n15_;
  assign new_n_n144_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n10_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n133_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n122_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n111_ = new_n_n27_ & new_n_n30_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n100_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n5_ = ~new_ns_;
  assign new_n_n894_ = new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n15_ & new_n_n24_ & new_n_n30_ & new_n_n18_ & new_n_n26_ & new_n_n25_ & new_n_n29_ & new_n_n16_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n885_ = new_n_n33_ & new_n_n34_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nk0_ & new_nd0_ & new_n_n23_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n872_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_ni0_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n863_ = new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_nk0_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n795_ = new_n_n4_ & new_n_n6_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n3_ & new_nk0_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n787_ = new_n_n25_ & new_n_n26_ & new_nv_ & new_n_n27_ & new_n_n24_ & new_nd0_ & new_nj0_ & new_n_n22_;
  assign new_n_n774_ = new_n_n22_ & new_n_n24_ & new_n_n25_ & new_n_n26_ & new_nz_ & new_nu_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nh0_;
  assign new_n_n765_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_nc_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n31_;
  assign new_n_n697_ = new_n_n20_ & new_n_n27_ & new_nl0_ & new_n_n14_ & new_n_n24_ & new_n_n22_ & new_nj0_ & new_nf0_ & new_n_n26_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n688_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nl0_ & new_n_n14_ & new_n_n26_ & new_n_n23_ & new_n_n24_ & new_n_n0_ & new_n_n34_ & new_n_n1_ & new_n_n33_ & new_n_n17_;
  assign new_n_n675_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_nl0_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n666_ = new_n_n31_ & new_n_n17_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n23_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n33_;
  assign new_n_n639_ = new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_n_n15_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n7_ & new_n_n21_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n598_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n576_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_ & new_n_n30_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n16_ & new_n_n5_ & new_nd_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n567_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n28_ & new_n_n31_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n22_ & new_n_n16_ & new_nj0_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n550_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_no_ & new_nh0_;
  assign new_n_n541_ = new_no_ & new_nn_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_ne0_;
  assign new_n_n478_ = new_nr_ & new_nm_ & new_n_n30_ & new_ng0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n469_ = new_n_n14_ & new_nm0_ & new_n_n20_ & new_n_n1_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_n_n24_;
  assign new_n_n451_ = new_n_n25_ & new_nm0_ & new_n_n10_ & new_n_n14_ & new_n_n20_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_n_n15_;
  assign new_n_n442_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n24_ & new_n_n1_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n420_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n2_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n379_ = new_n_n15_ & new_n_n26_ & new_n_n14_ & new_nm0_ & new_n_n10_ & new_n_n20_ & new_nt_ & new_n_n9_ & new_nj_ & new_n_n30_ & new_n_n34_ & new_n_n29_ & new_n_n27_;
  assign new_n_n352_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n343_ = new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_nt_ & new_n_n10_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n330_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n11_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n321_ = new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_n_n15_;
  assign new_n_n253_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n2_ & new_n_n22_ & new_n_n16_ & new_n_n27_ & new_n_n6_ & new_n_n24_ & new_nj0_;
  assign new_n_n244_ = new_n_n29_ & new_n_n8_ & new_nm0_ & new_n_n27_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n3_ & new_n_n10_ & new_n_n1_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n231_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n222_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_nd_ & new_n_n1_ & new_n_n11_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n200_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n10_ & new_n_n25_ & new_nk_ & new_nm_ & new_nt_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n8_;
  assign new_n_n154_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n25_ & new_nm0_ & new_n_n3_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n145_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n11_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n132_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n123_ = new_n_n29_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n110_ = new_n_n27_ & new_n_n8_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n101_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n7_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n6_ = ~new_nj_;
  assign new_n_n893_ = new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n15_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n25_ & new_n_n21_ & new_n_n16_ & new_n_n33_ & new_n_n10_ & new_n_n32_ & new_n_n31_;
  assign new_n_n882_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nj0_ & new_n_n22_ & new_n_n23_ & new_n_n21_ & new_n_n24_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n875_ = new_n_n34_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n864_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_ni0_ & new_n_n20_ & new_n_n21_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n848_ = new_n_n27_ & new_n_n28_ & new_n_n15_ & new_nd0_ & new_nk0_ & new_n_n18_ & new_n_n24_ & new_n_n25_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n33_ & new_n_n31_;
  assign new_n_n794_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n28_ & new_n_n31_ & new_nk0_ & new_n_n15_ & new_nd0_ & new_n_n27_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n784_ = new_n_n26_ & new_n_n22_ & new_nv_ & new_n_n25_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_nd0_ & new_n_n24_;
  assign new_n_n777_ = new_n_n28_ & new_n_n29_ & new_nh0_ & new_n_n27_ & new_nz_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n766_ = new_n_n21_ & new_nj0_ & new_n_n23_ & new_n_n22_ & new_nv_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nd0_;
  assign new_n_n750_ = new_n_n20_ & new_n_n27_ & new_n_n22_ & new_nj0_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n739_ = new_n_n27_ & new_n_n28_ & new_n_n21_ & new_nh0_ & new_ni0_ & new_nz_ & new_n_n33_ & new_nu_ & new_n_n32_ & new_n_n31_ & new_n_n30_;
  assign new_n_n696_ = new_n_n27_ & new_n_n28_ & new_n_n14_ & new_n_n20_ & new_nl0_ & new_n_n23_ & new_n_n24_ & new_nf0_ & new_n_n26_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n29_;
  assign new_n_n685_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n33_;
  assign new_n_n678_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_nl0_ & new_nj0_ & new_n_n24_ & new_n_n23_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n33_;
  assign new_n_n667_ = new_n_n17_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n15_ & new_nl0_ & new_nd0_ & new_n_n23_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n651_ = new_nn_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_nj0_ & new_nl0_ & new_n_n20_ & new_n_n22_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n640_ = new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_n_n24_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n7_ & new_n_n21_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n597_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n15_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n586_ = new_n_n33_ & new_n_n6_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n568_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nd_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n22_ & new_n_n16_ & new_nj0_ & new_n_n5_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n553_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ne0_ & new_nx_;
  assign new_n_n542_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_nf0_ & new_nb0_;
  assign new_n_n499_ = new_nu_ & new_n_n19_ & new_nj0_ & new_n_n27_ & new_nd0_ & new_n_n22_;
  assign new_n_n488_ = new_n_n22_ & new_no_ & new_nn_ & new_n_n27_ & new_nw_ & new_ng0_ & new_nj0_;
  assign new_n_n454_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n20_ & new_n_n30_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n26_;
  assign new_n_n443_ = new_n_n15_ & new_n_n26_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n410_ = new_n_n27_ & new_n_n8_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n20_ & new_nm0_ & new_ni0_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n30_;
  assign new_n_n389_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n24_ & new_n_n27_ & new_nj0_ & new_nm0_;
  assign new_n_n355_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_n_n22_ & new_n_n20_ & new_n_n23_ & new_n_n16_ & new_nj0_ & new_n_n27_ & new_nm0_ & new_n_n14_;
  assign new_n_n344_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_nt_ & new_n_n10_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n311_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n10_ & new_n_n14_ & new_n_n9_ & new_nt_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n300_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n10_ & new_nm0_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n19_ & new_n_n30_;
  assign new_n_n256_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n245_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n24_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n3_ & new_n_n1_ & new_n_n11_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n230_ = new_n_n24_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n212_ = new_nm0_ & new_n_n27_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n201_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n14_ & new_n_n25_ & new_nk_ & new_nm_ & new_nt_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n29_;
  assign new_n_n157_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n2_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n27_ & new_n_n24_;
  assign new_n_n146_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n11_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n131_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n120_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n113_ = new_n_n27_ & new_n_n30_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n102_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n7_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n7_ = ~new_nb_;
  assign new_n_n892_ = new_n_n15_ & new_n_n27_ & new_n_n24_ & new_nk0_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n25_ & new_n_n21_ & new_n_n16_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n883_ = new_n_n33_ & new_n_n10_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n22_ & new_n_n20_ & new_n_n23_ & new_n_n21_ & new_nk0_ & new_nj0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n874_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n24_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n865_ = new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_n_n30_ & new_nk0_ & new_ni0_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n838_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n30_ & new_n_n18_ & new_nk0_ & new_n_n15_ & new_n_n21_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n793_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n5_ & new_nd_ & new_nk0_ & new_nd0_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n785_ = new_n_n26_ & new_ni0_ & new_nv_ & new_n_n25_ & new_n_n31_ & new_n_n27_ & new_n_n30_ & new_nd0_ & new_n_n24_;
  assign new_n_n776_ = new_n_n27_ & new_n_n28_ & new_n_n23_ & new_nh0_ & new_nz_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n29_;
  assign new_n_n767_ = new_nj0_ & new_nd0_ & new_n_n23_ & new_n_n22_ & new_nv_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n749_ = new_nj0_ & new_n_n27_ & new_n_n22_ & new_n_n21_ & new_n_n23_ & new_nf0_ & new_nh_ & new_nu_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n740_ = new_n_n27_ & new_n_n28_ & new_nh0_ & new_n_n20_ & new_ni0_ & new_nz_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n695_ = new_n_n20_ & new_n_n27_ & new_nl0_ & new_n_n14_ & new_n_n24_ & new_n_n23_ & new_ni0_ & new_nf0_ & new_n_n26_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n28_;
  assign new_n_n686_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n14_ & new_n_n24_ & new_nl0_ & new_n_n26_ & new_n_n23_ & new_n_n15_ & new_n_n0_ & new_n_n33_ & new_n_n34_ & new_n_n17_ & new_n_n31_;
  assign new_n_n677_ = new_n_n31_ & new_n_n32_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_nl0_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n33_;
  assign new_n_n668_ = new_n_n17_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n24_ & new_nl0_ & new_nd0_ & new_n_n23_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n650_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_nj0_ & new_n_n24_ & new_nl0_ & new_n_n22_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n641_ = new_n_n33_ & new_n_n10_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n7_ & new_n_n21_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n596_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n34_;
  assign new_n_n587_ = new_n_n4_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n31_ & new_n_n17_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n21_ & new_n_n24_ & new_nl0_ & new_nd0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n578_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_nd_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n16_ & new_n_n15_ & new_n_n24_ & new_n_n5_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n34_;
  assign new_n_n552_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ng0_ & new_nx_;
  assign new_n_n543_ = new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ng0_ & new_nb0_;
  assign new_n_n498_ = new_nv_ & new_n_n19_ & new_n_n27_ & new_n_n30_ & new_nd0_ & new_ni0_;
  assign new_n_n489_ = new_n_n22_ & new_no_ & new_nn_ & new_n_n27_ & new_nw_ & new_ne0_ & new_nj0_;
  assign new_n_n453_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n20_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_n_n24_;
  assign new_n_n444_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n10_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n400_ = new_nm0_ & new_n_n27_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n7_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n399_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n7_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n354_ = new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n345_ = new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_nt_ & new_n_n14_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n310_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_n_n15_ & new_n_n24_ & new_nm_ & new_nm0_ & new_nj_ & new_n_n34_ & new_nl_ & new_ns_ & new_n_n19_;
  assign new_n_n301_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n19_ & new_n_n30_;
  assign new_n_n255_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n27_ & new_nm0_;
  assign new_n_n246_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n3_ & new_n_n1_ & new_n_n11_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n220_ = new_n_n29_ & new_n_n8_ & new_nm0_ & new_n_n27_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_nd_ & new_n_n10_ & new_n_n1_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n211_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n202_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n25_ & new_nm0_ & new_nk_ & new_nm_ & new_nt_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n8_;
  assign new_n_n156_ = new_nm0_ & new_n_n15_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n27_;
  assign new_n_n147_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_n_n3_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n130_ = new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_nm0_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n121_ = new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n112_ = new_n_n8_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n103_ = new_n_n29_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n7_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n8_ = ~new_nz_;
  assign new_n_n891_ = new_n_n34_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n23_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n880_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nk0_ & new_ni0_ & new_n_n23_ & new_n_n21_ & new_n_n30_ & new_n_n24_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n869_ = new_n_n34_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_nk0_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n858_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n15_ & new_ni0_ & new_n_n25_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n34_;
  assign new_n_n828_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n15_ & new_n_n2_ & new_n_n29_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n792_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n5_ & new_nd_ & new_nk0_ & new_n_n15_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n782_ = new_n_n28_ & new_n_n29_ & new_n_n21_ & new_n_n27_ & new_nf0_ & new_nh_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n771_ = new_nd0_ & new_n_n27_ & new_n_n22_ & new_nj0_ & new_nv_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n760_ = new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n20_ & new_ni0_ & new_nf0_ & new_nh_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n730_ = new_nj0_ & new_nh0_ & new_n_n22_ & new_n_n21_ & new_n_n23_ & new_nz_ & new_n_n33_ & new_n_n31_ & new_nu_ & new_n_n28_ & new_n_n27_;
  assign new_n_n719_ = new_nl0_ & new_n_n20_ & new_nj0_ & new_n_n24_ & new_n_n21_ & new_n_n26_ & new_n_n22_ & new_nf0_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n27_;
  assign new_n_n694_ = new_n_n14_ & new_n_n20_ & new_n_n24_ & new_nl0_ & new_nj0_ & new_n_n23_ & new_n_n22_ & new_nf0_ & new_n_n26_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n683_ = new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n672_ = new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n24_ & new_nl0_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n33_ & new_n_n32_;
  assign new_n_n661_ = new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_n_n14_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n15_ & new_nl0_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n34_;
  assign new_n_n631_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_nj0_ & new_nl0_ & new_n_n14_ & new_n_n7_ & new_n_n22_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n620_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n5_ & new_nd_ & new_nl0_ & new_n_n20_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n609_ = new_n_n4_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n28_ & new_n_n31_ & new_nj0_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n595_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nj0_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n2_ & new_n_n22_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n584_ = new_n_n33_ & new_n_n6_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n21_ & new_n_n15_ & new_n_n5_ & new_nd_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n573_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n30_ & new_n_n31_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n16_ & new_n_n15_ & new_nl0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n562_ = new_n_n33_ & new_n_n34_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n2_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n533_ = new_n_n22_ & new_nw_ & new_nj0_ & new_n_n27_ & new_no_ & new_nh0_;
  assign new_n_n522_ = new_nq_ & new_nw_ & new_ne0_ & new_n_n27_ & new_nj0_ & new_n_n22_;
  assign new_n_n511_ = new_nb0_ & new_n_n30_ & new_ng0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n500_ = new_nu_ & new_n_n19_ & new_n_n27_ & new_n_n30_ & new_nd0_ & new_ni0_;
  assign new_n_n497_ = new_nv_ & new_n_n19_ & new_nj0_ & new_n_n27_ & new_nd0_ & new_n_n22_;
  assign new_n_n486_ = new_n_n22_ & new_n_n20_ & new_nn_ & new_ne0_ & new_n_n27_ & new_nj0_ & new_no_;
  assign new_n_n475_ = new_nr_ & new_nm_ & new_nw_ & new_ng0_ & new_n_n27_ & new_nj0_ & new_n_n22_;
  assign new_n_n464_ = new_n_n10_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n27_ & new_n_n8_ & new_n_n26_ & new_nm0_;
  assign new_n_n434_ = new_n_n15_ & new_n_n24_ & new_n_n20_ & new_nm0_ & new_ni0_ & new_n_n2_ & new_nj_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n26_;
  assign new_n_n423_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n2_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n412_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_nt_ & new_n_n10_ & new_n_n20_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n401_ = new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n398_ = new_nm0_ & new_n_n24_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n7_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n387_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_n_n22_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_nj0_ & new_n_n27_ & new_nm0_ & new_n_n14_;
  assign new_n_n376_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n10_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n8_;
  assign new_n_n365_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n23_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n335_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n324_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n25_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n313_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n9_ & new_nt_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n302_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n19_ & new_n_n30_;
  assign new_n_n299_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n10_ & new_n_n14_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n19_ & new_n_n30_;
  assign new_n_n288_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n25_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n277_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n24_ & new_n_n14_ & new_nt_ & new_n_n1_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n29_;
  assign new_n_n266_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n2_ & new_n_n1_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n250_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n25_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n236_ = new_n_n27_ & new_n_n29_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n20_ & new_n_n3_ & new_n_n10_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n225_ = new_nm0_ & new_nj0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n22_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n27_ & new_n_n24_;
  assign new_n_n214_ = new_n_n24_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n203_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n14_ & new_n_n25_ & new_nk_ & new_nm_ & new_n_n10_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n189_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n13_ & new_n_n14_ & new_n_n2_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n178_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n7_ & new_n_n11_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n167_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n27_ & new_n_n15_;
  assign new_n_n151_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n13_ & new_n_n14_ & new_n_n3_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n140_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n25_ & new_nd_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n137_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n13_ & new_n_n14_ & new_nd_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n126_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n115_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n104_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n7_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n79_ = new_n_n30_ & new_n_n19_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n68_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n1_ = ~new_nh_;
  assign new_n_n890_ = new_n_n33_ & new_n_n34_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n22_ & new_n_n20_ & new_n_n23_ & new_n_n24_ & new_nk0_ & new_nj0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n881_ = new_n_n33_ & new_n_n10_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_ni0_ & new_n_n20_ & new_n_n23_ & new_n_n21_ & new_n_n30_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n868_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nk0_ & new_n_n27_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n24_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n859_ = new_n_n33_ & new_n_n34_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_ni0_ & new_n_n20_ & new_n_n25_ & new_n_n30_ & new_nk0_ & new_n_n15_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n818_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nk0_ & new_n_n15_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n24_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n34_;
  assign new_n_n791_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n28_ & new_n_n31_ & new_n_n24_ & new_nk0_ & new_nd0_ & new_n_n27_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n783_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n770_ = new_nj0_ & new_nd0_ & new_n_n22_ & new_n_n21_ & new_nv_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n27_;
  assign new_n_n761_ = new_n_n28_ & new_n_n30_ & new_n_n21_ & new_n_n27_ & new_ni0_ & new_nf0_ & new_nh_ & new_n_n32_ & new_n_n33_ & new_nu_ & new_n_n31_;
  assign new_n_n729_ = new_n_n28_ & new_n_n29_ & new_n_n20_ & new_n_n27_ & new_nl0_ & new_n_n21_ & new_n_n15_ & new_n_n26_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n720_ = new_n_n20_ & new_n_n27_ & new_n_n24_ & new_nl0_ & new_n_n21_ & new_n_n26_ & new_ni0_ & new_nf0_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n28_;
  assign new_n_n693_ = new_n_n17_ & new_n_n32_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n26_ & new_nl0_ & new_n_n14_ & new_n_n0_ & new_n_n10_ & new_n_n1_ & new_n_n34_ & new_n_n33_;
  assign new_n_n684_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n24_ & new_nl0_ & new_n_n23_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n33_ & new_n_n31_;
  assign new_n_n671_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_n_n22_ & new_n_n16_ & new_n_n21_ & new_nj0_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n662_ = new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_n_n14_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n24_ & new_nl0_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n34_;
  assign new_n_n630_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n14_ & new_n_n20_ & new_n_n16_ & new_nj0_ & new_n_n24_ & new_nl0_ & new_n_n7_ & new_n_n22_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n34_;
  assign new_n_n621_ = new_n_n33_ & new_n_n4_ & new_n_n3_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n599_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_ & new_n_n30_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n2_ & new_ni0_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n594_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_n_n2_ & new_n_n22_ & new_n_n16_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n585_ = new_n_n4_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n31_ & new_n_n17_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n21_ & new_n_n15_ & new_nl0_ & new_nd0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n572_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nd_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n15_ & new_n_n5_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n563_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n2_ & new_n_n15_ & new_nl0_ & new_n_n14_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n532_ = new_n_n22_ & new_n_n27_ & new_nj0_ & new_ne0_ & new_nx_ & new_n_n20_;
  assign new_n_n523_ = new_nq_ & new_n_n30_ & new_nf0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n510_ = new_nb0_ & new_n_n30_ & new_nf0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n501_ = new_nr_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_nf0_ & new_nm_;
  assign new_n_n496_ = new_nd0_ & new_no_ & new_nn_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n487_ = new_n_n22_ & new_no_ & new_nn_ & new_n_n27_ & new_nw_ & new_nj0_ & new_nf0_;
  assign new_n_n474_ = new_nr_ & new_nm_ & new_nw_ & new_nj0_ & new_n_n27_ & new_nf0_ & new_n_n22_;
  assign new_n_n465_ = new_n_n1_ & new_n_n14_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_;
  assign new_n_n433_ = new_nm0_ & new_n_n15_ & new_n_n20_ & new_n_n14_ & new_ni0_ & new_n_n2_ & new_nj_ & new_n_n27_ & new_n_n30_ & new_n_n26_ & new_n_n24_;
  assign new_n_n424_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n2_ & new_n_n10_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n411_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_nt_ & new_n_n10_ & new_n_n20_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n402_ = new_n_n24_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n397_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n7_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n388_ = new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n10_ & new_n_n22_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n27_ & new_n_n8_ & new_nj0_ & new_nm0_;
  assign new_n_n375_ = new_n_n15_ & new_n_n26_ & new_n_n14_ & new_nm0_ & new_n_n10_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n27_;
  assign new_n_n366_ = new_nm0_ & new_n_n24_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n1_ & new_n_n23_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n334_ = new_nj0_ & new_n_n24_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n325_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n312_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n10_ & new_nm0_ & new_n_n9_ & new_nt_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n303_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_n_n10_ & new_n_n14_ & new_nm_ & new_nt_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n298_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_nt_ & new_nm0_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n289_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n276_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n26_ & new_n_n1_ & new_nt_ & new_n_n10_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n8_;
  assign new_n_n267_ = new_nm0_ & new_n_n26_ & new_n_n1_ & new_n_n14_ & new_n_n10_ & new_n_n9_ & new_nt_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n240_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n235_ = new_nm0_ & new_n_n27_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n20_ & new_n_n3_ & new_n_n10_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n226_ = new_nj0_ & new_n_n24_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n22_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n213_ = new_nm0_ & new_n_n24_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n204_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n25_ & new_nm0_ & new_nk_ & new_nm_ & new_n_n10_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n199_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n10_ & new_n_n14_ & new_nk_ & new_nm_ & new_nt_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n29_;
  assign new_n_n177_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n7_ & new_n_n11_ & new_n_n16_ & new_n_n19_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_n_n168_ = new_nm0_ & new_n_n15_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n8_ & new_n_n27_;
  assign new_n_n150_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n25_ & new_n_n20_ & new_n_n3_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n141_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n14_ & new_n_n25_ & new_nd_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n136_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_nd_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n127_ = new_n_n30_ & new_n_n19_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n114_ = new_n_n8_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n105_ = new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n7_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n78_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n69_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n2_ = ~new_nk_;
  assign new_n_n889_ = new_n_n34_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n23_ & new_n_n30_ & new_nk0_ & new_ni0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n878_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n24_ & new_nk0_ & new_n_n23_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n871_ = new_n_n34_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_nk0_ & new_n_n20_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n860_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n24_ & new_nk0_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n808_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n20_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n790_ = new_n_n33_ & new_n_n34_ & new_n_n3_ & new_n_n32_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nk0_ & new_n_n15_ & new_nd0_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n4_;
  assign new_n_n780_ = new_n_n27_ & new_n_n28_ & new_n_n23_ & new_n_n21_ & new_nf0_ & new_nh_ & new_n_n31_ & new_n_n33_ & new_n_n30_ & new_n_n29_;
  assign new_n_n773_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_nd0_ & new_nv_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n762_ = new_n_n28_ & new_n_n30_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n710_ = new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nl0_ & new_n_n14_ & new_n_n26_ & new_ni0_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n32_;
  assign new_n_n699_ = new_n_n28_ & new_n_n29_ & new_n_n20_ & new_n_n27_ & new_n_n14_ & new_n_n24_ & new_nl0_ & new_nf0_ & new_n_n26_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_n_n692_ = new_n_n31_ & new_n_n17_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n14_ & new_n_n27_ & new_n_n26_ & new_n_n24_ & new_nl0_ & new_n_n0_ & new_n_n34_ & new_n_n1_ & new_n_n33_ & new_n_n32_;
  assign new_n_n681_ = new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n15_ & new_nl0_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n33_;
  assign new_n_n674_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n24_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n33_;
  assign new_n_n663_ = new_n_n33_ & new_n_n34_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_ni0_ & new_n_n16_ & new_nl0_ & new_n_n14_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n629_ = new_n_n34_ & new_n_n10_ & new_n_n17_ & new_n_n33_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n23_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n611_ = new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n3_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n4_;
  assign new_n_n600_ = new_n_n32_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n29_ & new_n_n27_ & new_n_n28_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n2_ & new_n_n16_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n34_;
  assign new_n_n593_ = new_n_n34_ & new_n_n10_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n7_ & new_nl0_ & new_n_n14_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n582_ = new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n17_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_nd_ & new_nl0_ & new_nd0_ & new_n_n27_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_n_n5_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n575_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n30_ & new_n_n31_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n16_ & new_n_n24_ & new_nl0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n564_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n2_ & new_n_n24_ & new_nl0_ & new_n_n14_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n531_ = new_n_n22_ & new_n_n27_ & new_nj0_ & new_ng0_ & new_nx_ & new_n_n20_;
  assign new_n_n520_ = new_nq_ & new_nw_ & new_nj0_ & new_n_n27_ & new_nf0_ & new_n_n22_;
  assign new_n_n513_ = new_nb0_ & new_nw_ & new_n_n27_ & new_n_n30_ & new_nf0_ & new_ni0_;
  assign new_n_n502_ = new_nr_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ng0_ & new_nm_;
  assign new_n_n495_ = new_ni0_ & new_no_ & new_nn_ & new_n_n30_ & new_nw_ & new_n_n27_ & new_ne0_;
  assign new_n_n484_ = new_n_n22_ & new_n_n20_ & new_nn_ & new_nj0_ & new_n_n27_ & new_nf0_ & new_no_;
  assign new_n_n477_ = new_nr_ & new_nm_ & new_n_n30_ & new_nf0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n466_ = new_n_n1_ & new_nm0_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n27_ & new_n_n8_ & new_n_n26_ & new_n_n24_;
  assign new_n_n450_ = new_nm0_ & new_n_n15_ & new_n_n20_ & new_n_n25_ & new_ni0_ & new_n_n30_ & new_n_n27_ & new_n_n8_ & new_n_n26_ & new_n_n24_;
  assign new_n_n432_ = new_nm0_ & new_n_n15_ & new_n_n20_ & new_n_n10_ & new_ni0_ & new_n_n2_ & new_nj_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n26_;
  assign new_n_n421_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n2_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n414_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_nt_ & new_nm0_ & new_n_n20_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n403_ = new_n_n15_ & new_n_n26_ & new_n_n14_ & new_nm0_ & new_n_n10_ & new_n_n20_ & new_nt_ & new_ni0_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n27_;
  assign new_n_n396_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n7_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n29_ & new_n_n27_;
  assign new_n_n385_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n20_ & new_n_n14_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n29_;
  assign new_n_n378_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n8_;
  assign new_n_n367_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n23_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n351_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n24_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n1_ & new_n_n11_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n340_ = new_n_n27_ & new_n_n29_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n333_ = new_nm0_ & new_nj0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n27_ & new_n_n24_;
  assign new_n_n322_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n25_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n315_ = new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n9_ & new_n_n10_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n304_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n10_ & new_nm0_ & new_nm_ & new_nt_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n297_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_nt_ & new_n_n14_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n286_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n25_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n24_;
  assign new_n_n279_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n26_ & new_n_n14_ & new_n_n10_ & new_n_n1_ & new_nk_ & new_nm_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n268_ = new_n_n26_ & new_n_n27_ & new_n_n1_ & new_nm0_ & new_n_n10_ & new_n_n9_ & new_nt_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n252_ = new_n_n13_ & new_nm0_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_n_n22_ & new_n_n16_ & new_n_n8_ & new_n_n6_ & new_n_n27_ & new_nj0_;
  assign new_n_n241_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n13_ & new_n_n14_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n234_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n223_ = new_n_n14_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n27_ & new_nj0_;
  assign new_n_n216_ = new_n_n27_ & new_n_n29_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_nd_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n205_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n25_ & new_nm0_ & new_nk_ & new_nm_ & new_n_n14_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n198_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n25_ & new_nm0_ & new_nk_ & new_nm_ & new_n_n9_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n187_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n169_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n20_ & new_n_n11_ & new_n_n2_ & new_n_n7_ & new_ni0_ & new_n_n16_ & new_n_n30_ & new_nj_ & new_n_n27_ & new_n_n24_;
  assign new_n_n153_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n14_ & new_n_n25_ & new_n_n3_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n142_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n25_ & new_nm0_ & new_nd_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n135_ = new_n_n15_ & new_n_n27_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_nd_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n124_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n117_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n106_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n7_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n99_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n88_ = new_n_n27_ & new_n_n8_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n3_ = ~new_nt_;
  assign new_n_n888_ = new_n_n33_ & new_n_n34_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_ni0_ & new_n_n20_ & new_n_n23_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n879_ = new_n_n33_ & new_n_n10_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nk0_ & new_n_n20_ & new_n_n23_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n870_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_nk0_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n861_ = new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nk0_ & new_n_n27_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n798_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_nd_ & new_nk0_ & new_n_n15_ & new_n_n20_ & new_n_n29_ & new_n_n30_ & new_n_n5_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n789_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_nk0_ & new_n_n29_ & new_n_n30_ & new_n_n18_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n781_ = new_n_n28_ & new_n_n29_ & new_n_n23_ & new_n_n27_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n30_;
  assign new_n_n772_ = new_nd0_ & new_n_n27_ & new_ni0_ & new_n_n21_ & new_nv_ & new_n_n33_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n28_;
  assign new_n_n763_ = new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_ni0_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_nu_;
  assign new_n_n709_ = new_n_n28_ & new_n_n30_ & new_n_n20_ & new_n_n27_ & new_n_n14_ & new_n_n15_ & new_nl0_ & new_n_n26_ & new_ni0_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n700_ = new_n_n27_ & new_n_n28_ & new_n_n14_ & new_n_n20_ & new_nl0_ & new_n_n22_ & new_nj0_ & new_n_n26_ & new_n_n23_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n31_;
  assign new_n_n691_ = new_n_n31_ & new_n_n17_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_n_n14_ & new_n_n27_ & new_n_n26_ & new_n_n15_ & new_nl0_ & new_n_n0_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n32_;
  assign new_n_n682_ = new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_n_n24_ & new_nl0_ & new_n_n23_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n33_;
  assign new_n_n673_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n7_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n33_;
  assign new_n_n664_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_n_n14_ & new_n_n20_ & new_n_n16_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n23_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n34_ & new_n_n33_;
  assign new_n_n619_ = new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n3_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_n_n24_ & new_nl0_ & new_n_n20_ & new_n_n27_ & new_n_n16_ & new_n_n21_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n4_;
  assign new_n_n610_ = new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n30_ & new_n_n27_ & new_nl0_ & new_n_n20_ & new_n_n15_ & new_n_n24_ & new_n_n5_ & new_nd_ & new_ni0_ & new_n_n16_ & new_n_n21_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n6_ & new_n_n33_;
  assign new_n_n601_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n28_ & new_n_n29_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_n_n27_ & new_n_n2_ & new_n_n16_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n10_ & new_n_n6_;
  assign new_n_n592_ = new_n_n33_ & new_n_n34_ & new_n_n17_ & new_n_n32_ & new_n_n31_ & new_n_n29_ & new_n_n30_ & new_n_n14_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n7_ & new_n_n24_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n583_ = new_n_n33_ & new_n_n4_ & new_n_n3_ & new_n_n32_ & new_n_n17_ & new_n_n30_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n21_ & new_n_n15_ & new_n_n24_ & new_nl0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_n_n574_ = new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n32_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nd_ & new_nl0_ & new_n_n14_ & new_n_n20_ & new_ni0_ & new_n_n16_ & new_n_n24_ & new_n_n5_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n565_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_ & new_n_n17_ & new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n2_ & new_nl0_ & new_n_n14_ & new_nd0_ & new_n_n0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n530_ = new_n_n22_ & new_n_n27_ & new_nx_ & new_nj0_ & new_nf0_ & new_n_n20_;
  assign new_n_n521_ = new_nq_ & new_nw_ & new_ng0_ & new_n_n27_ & new_nj0_ & new_n_n22_;
  assign new_n_n512_ = new_nb0_ & new_n_n30_ & new_ne0_ & new_n_n27_ & new_n_n20_ & new_ni0_;
  assign new_n_n503_ = new_nr_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_ne0_ & new_nm_;
  assign new_n_n494_ = new_ni0_ & new_no_ & new_nn_ & new_n_n30_ & new_nw_ & new_n_n27_ & new_ng0_;
  assign new_n_n485_ = new_n_n22_ & new_n_n20_ & new_nn_ & new_ng0_ & new_n_n27_ & new_nj0_ & new_no_;
  assign new_n_n476_ = new_nr_ & new_nm_ & new_nw_ & new_ne0_ & new_n_n27_ & new_nj0_ & new_n_n22_;
  assign new_n_n467_ = new_n_n1_ & new_n_n14_ & new_n_n20_ & new_n_n10_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n26_ & new_nm0_;
  assign new_n_n440_ = new_n_n26_ & new_n_n27_ & new_n_n1_ & new_nm0_ & new_n_n10_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n431_ = new_n_n14_ & new_nm0_ & new_n_n20_ & new_n_n10_ & new_ni0_ & new_n_n2_ & new_nj_ & new_n_n27_ & new_n_n30_ & new_n_n26_ & new_n_n15_;
  assign new_n_n422_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n2_ & new_nm_ & new_nj_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n413_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_nt_ & new_n_n14_ & new_n_n20_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n404_ = new_n_n26_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n10_ & new_n_n20_ & new_nt_ & new_ni0_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n395_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n7_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nm0_;
  assign new_n_n386_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n20_ & new_nm0_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n8_;
  assign new_n_n377_ = new_n_n24_ & new_n_n26_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_ni0_ & new_n_n20_ & new_n_n9_ & new_nj_ & new_n_n34_ & new_nl_ & new_n_n30_ & new_n_n27_;
  assign new_n_n368_ = new_nm0_ & new_n_n27_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n23_ & new_n_n16_ & new_n_n30_ & new_n_n19_ & new_n_n8_ & new_n_n29_;
  assign new_n_n350_ = new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n8_ & new_n_n27_ & new_n_n15_ & new_n_n26_ & new_n_n10_ & new_nm0_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_ns_;
  assign new_n_n341_ = new_n_n24_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n20_ & new_n_n1_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n332_ = new_nm0_ & new_nj0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n323_ = new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_n_n20_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n15_;
  assign new_n_n314_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n9_ & new_nt_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n305_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_nm_ & new_nt_ & new_nj_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n296_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n26_ & new_nm0_ & new_nt_ & new_n_n10_ & new_nm_ & new_n_n9_ & new_nj_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n8_;
  assign new_n_n287_ = new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n20_ & new_n_n16_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n15_;
  assign new_n_n278_ = new_n_n27_ & new_n_n29_ & new_n_n24_ & new_n_n26_ & new_nm0_ & new_nt_ & new_n_n1_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n19_ & new_ns_ & new_n_n30_ & new_n_n8_;
  assign new_n_n269_ = new_n_n24_ & new_n_n26_ & new_n_n14_ & new_nm0_ & new_n_n1_ & new_n_n9_ & new_nt_ & new_nk_ & new_nm_ & new_n_n34_ & new_n_n30_ & new_n_n19_ & new_n_n29_ & new_n_n27_;
  assign new_n_n251_ = new_n_n13_ & new_n_n14_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n20_ & new_n_n10_ & new_n_n2_ & new_n_n22_ & new_n_n16_ & new_n_n27_ & new_n_n6_ & new_nj0_ & new_nm0_;
  assign new_n_n242_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n25_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n233_ = new_n_n15_ & new_n_n24_ & new_n_n25_ & new_nm0_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n16_ & new_nn_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n224_ = new_nm0_ & new_nj0_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_ & new_n_n1_ & new_n_n22_ & new_n_n20_ & new_n_n3_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n8_ & new_n_n27_;
  assign new_n_n215_ = new_nm0_ & new_n_n27_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n1_ & new_n_n11_ & new_nd_ & new_n_n20_ & new_n_n10_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n29_;
  assign new_n_n206_ = new_n_n29_ & new_n_n8_ & new_n_n26_ & new_n_n27_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_nk_ & new_nm_ & new_n_n25_ & new_nl_ & new_ns_ & new_n_n34_ & new_n_n19_ & new_n_n30_;
  assign new_n_n197_ = new_n_n26_ & new_n_n27_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n14_ & new_n_n25_ & new_nk_ & new_nm_ & new_n_n9_ & new_nl_ & new_n_n19_ & new_n_n34_ & new_n_n30_ & new_n_n29_;
  assign new_n_n188_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_n_n2_ & new_n_n10_ & new_n_n11_ & new_n_n16_ & new_n_n19_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n179_ = new_n_n25_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n2_ & new_ni0_ & new_n_n20_ & new_n_n16_ & new_n_n30_ & new_n_n6_ & new_n_n27_ & new_n_n15_;
  assign new_n_n152_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n25_ & new_n_n3_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n19_ & new_n_n30_;
  assign new_n_n143_ = new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n25_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_n_n3_ & new_n_n10_ & new_n_n16_ & new_n_n4_ & new_n_n6_ & new_n_n30_ & new_n_n27_;
  assign new_n_n134_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n25_ & new_n_n12_ & new_n_n13_ & new_nd_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n16_ & new_n_n5_ & new_n_n6_ & new_n_n30_ & new_n_n8_;
  assign new_n_n125_ = new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n19_;
  assign new_n_n116_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n107_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n7_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_n_n98_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n7_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n89_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n7_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n9_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n4_ = ~new_nl_;
  assign new_n_n54_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n9_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n43_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_ny0_ = new_n_n27_ & new_n_n28_ & new_nh0_ & new_n_n20_ & new_n_n22_ & new_nj0_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_n_n31_ & new_nz_;
  assign new_nj1_ = new_n_n28_ & new_nz_ & new_n_n20_ & new_n_n27_ & new_nh0_ & new_ni0_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_n_n31_ & new_n_n30_;
  assign new_nu1_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nd0_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_nv_ & new_n_n19_;
  assign new_n_n55_ = new_n_n29_ & new_n_n30_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n9_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n42_ = new_n_n27_ & new_n_n8_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_nx0_ = new_n_n31_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_nc_ & new_n_n34_ & new_n_n23_ & new_n_n33_ & new_n_n17_;
  assign new_nk1_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_nd0_ & new_nj0_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_nw_ & new_n_n31_;
  assign new_nt1_ = new_n_n28_ & new_n_n30_ & new_n_n20_ & new_n_n27_ & new_nh0_ & new_ni0_ & new_n_n23_ & new_no_ & new_n_n34_ & new_n_n33_ & new_n_n31_;
  assign new_n_n56_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n9_ & new_n_n10_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n41_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_na1_ = new_n_n31_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_nu_ & new_n_n18_;
  assign new_nh1_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_nd0_ & new_nj0_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_nw_ & new_n_n31_;
  assign new_ns1_ = new_nh0_ & new_n_n24_ & new_nj0_ & new_n_n22_ & new_no_ & new_n_n20_ & new_n_n27_ & new_n_n26_ & new_n_n25_;
  assign new_n_n57_ = new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n14_ & new_nm0_ & new_n_n9_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_n_n40_ = new_n_n27_ & new_n_n8_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_nz0_ = new_n_n27_ & new_n_n28_ & new_nh0_ & new_n_n20_ & new_n_n22_ & new_nj0_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_nz_;
  assign new_ni1_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_nd0_ & new_nj0_ & new_n_n23_ & new_n_n33_ & new_n_n34_ & new_nw_ & new_n_n31_;
  assign new_nr1_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nd0_ & new_n_n23_ & new_n_n33_ & new_n_n34_ & new_nv_ & new_n_n19_;
  assign new_n_n0_ = ~new_na_;
  assign new_n_n877_ = new_n_n31_ & new_n_n33_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_n_n18_ & new_nk0_ & new_n_n23_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n866_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n22_ & new_n_n20_ & new_n_n21_ & new_n_n24_ & new_nk0_ & new_nj0_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n768_ = new_n_n21_ & new_nd0_ & new_n_n23_ & new_ni0_ & new_nv_ & new_n_n33_ & new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n27_;
  assign new_n_n58_ = new_n_n8_ & new_n_n30_ & new_n_n27_ & new_n_n29_ & new_n_n24_ & new_nm0_ & new_n_n15_ & new_n_n9_ & new_n_n11_ & new_n_n12_ & new_n_n13_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n19_;
  assign new_nb2_ = new_n_n22_ & new_n_n24_ & new_nj0_ & new_nw_ & new_nd0_ & new_n_n27_ & new_n_n26_ & new_n_n25_;
  assign new_n_n32_ = ~new_nr_;
  assign new_n_n21_ = ~new_no_;
  assign new_n_n10_ = ~new_ni_;
  assign new_n_n876_ = new_n_n28_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_nk0_ & new_n_n18_ & new_n_n24_ & new_n_n23_ & new_n_n21_ & new_n_n29_ & new_n_n30_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n33_;
  assign new_n_n867_ = new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_nk0_ & new_nj0_ & new_n_n22_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n778_ = new_n_n21_ & new_nj0_ & new_n_n26_ & new_n_n22_ & new_n_n25_ & new_n_n1_ & new_n_n20_ & new_n_n27_ & new_nl0_ & new_n_n24_;
  assign new_n_n59_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_ns_ & new_n_n30_;
  assign new_nc2_ = new_n_n28_ & new_n_n30_ & new_nd0_ & new_n_n27_ & new_ni0_ & new_n_n23_ & new_n_n33_ & new_n_n34_ & new_nw_ & new_n_n31_;
  assign new_n_n33_ = ~new_nq_;
  assign new_n_n20_ = ~new_nd0_;
  assign new_n_n11_ = ~new_ng_;
  assign new_n_n897_ = new_nk0_ & new_n_n15_ & new_n_n30_ & new_n_n18_ & new_n_n29_ & new_n_n25_ & new_n_n21_ & new_n_n26_ & new_n_n23_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n886_ = new_n_n33_ & new_n_n34_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nk0_ & new_n_n20_ & new_n_n23_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_no0_ = new_n_n668_ | new_ni1_ | new_n_n650_ | new_n_n659_ | new_n_n632_ | new_n_n641_ | new_n_n598_ | new_n_n623_ | new_n_n580_ | new_n_n589_ | new_n_n562_ | new_n_n571_ | new_n_n669_ | new_nh1_ | new_n_n651_ | new_n_n658_ | new_n_n633_ | new_n_n640_ | new_n_n608_ | new_n_n622_ | new_n_n579_ | new_n_n590_ | new_n_n561_ | new_n_n572_ | new_nk1_ | new_n_n554_ | new_n_n679_ | new_n_n688_ | new_n_n643_ | new_n_n652_ | new_n_n630_ | new_n_n591_ | new_n_n621_ | new_n_n569_ | new_n_n582_ | new_n_n555_ | new_n_n560_ | new_n_n689_ | new_nj1_ | new_n_n653_ | new_n_n678_ | new_n_n631_ | new_n_n642_ | new_n_n592_ | new_n_n620_ | new_n_n570_ | new_n_n581_ | new_n_n556_ | new_n_n559_ | new_n_n681_ | new_n_n690_ | new_n_n663_ | new_n_n672_ | new_n_n619_ | new_n_n628_ | new_n_n584_ | new_n_n593_ | new_n_n566_ | new_n_n575_ | new_n_n691_ | new_nl1_ | new_n_n673_ | new_n_n680_ | new_n_n662_ | new_n_n618_ | new_n_n629_ | new_n_n583_ | new_n_n594_ | new_n_n565_ | new_n_n576_ | new_n_n683_ | new_n_n692_ | new_n_n661_ | new_n_n670_ | new_n_n639_ | new_n_n648_ | new_n_n586_ | new_n_n595_ | new_n_n564_ | new_n_n573_ | new_n_n682_ | new_n_n693_ | new_n_n660_ | new_n_n671_ | new_n_n638_ | new_n_n649_ | new_n_n585_ | new_n_n596_ | new_n_n563_ | new_n_n574_ | new_n_n749_ | new_n_n758_ | new_n_n731_ | new_n_n740_ | new_n_n694_ | new_n_n722_ | new_n_n685_ | new_n_n667_ | new_n_n676_ | new_n_n759_ | new_n_n597_ | new_n_n741_ | new_n_n748_ | new_n_n723_ | new_n_n730_ | new_n_n684_ | new_n_n695_ | new_n_n666_ | new_n_n677_ | new_n_n760_ | new_n_n587_ | new_n_n738_ | new_n_n751_ | new_n_n724_ | new_n_n729_ | new_n_n687_ | new_n_n696_ | new_n_n665_ | new_n_n674_ | new_n_n761_ | new_n_n577_ | new_n_n739_ | new_n_n750_ | new_n_n725_ | new_n_n728_ | new_n_n686_ | new_n_n697_ | new_n_n664_ | new_n_n675_ | new_n_n567_ | new_na2_ | new_nn1_ | new_n_n753_ | new_n_n762_ | new_n_n735_ | new_n_n744_ | new_n_n654_ | new_n_n718_ | new_n_n636_ | new_n_n645_ | new_n_n557_ | new_n_n627_ | new_nb2_ | new_nm1_ | new_n_n752_ | new_n_n763_ | new_n_n734_ | new_n_n745_ | new_n_n655_ | new_n_n719_ | new_n_n637_ | new_n_n644_ | new_n_n786_ | new_n_n626_ | new_n_n764_ | new_n_n777_ | new_n_n742_ | new_n_n755_ | new_n_n720_ | new_n_n733_ | new_n_n647_ | new_n_n656_ | new_n_n634_ | new_n_n787_ | new_n_n625_ | new_n_n765_ | new_n_n776_ | new_n_n743_ | new_n_n754_ | new_n_n721_ | new_n_n732_ | new_n_n646_ | new_n_n657_ | new_n_n624_ | new_n_n635_ | new_ne2_ | new_nr1_ | new_n_n775_ | new_n_n784_ | new_n_n757_ | new_n_n766_ | new_nf2_ | new_nq1_ | new_n_n774_ | new_n_n785_ | new_n_n756_ | new_n_n767_ | new_nc2_ | new_np1_ | new_n_n773_ | new_n_n782_ | new_n_n737_ | new_n_n746_ | new_nd2_ | new_no1_ | new_n_n783_ | new_n_n747_ | new_n_n772_ | new_ny1_ | new_n_n736_ | new_n_n780_ | new_ni2_ | new_n_n726_ | new_n_n771_ | new_n_n707_ | new_n_n716_ | new_nj2_ | new_nx1_ | new_n_n770_ | new_n_n781_ | new_n_n717_ | new_n_n727_ | new_nw1_ | new_n_n706_ | new_n_n778_ | new_ng2_ | new_n_n714_ | new_n_n769_ | new_n_n617_ | new_n_n705_ | new_nh2_ | new_nu1_ | new_n_n768_ | new_n_n779_ | new_n_n704_ | new_n_n715_ | new_n_n712_ | new_n_n607_ | new_n_n703_ | new_n_n606_ | new_n_n615_ | new_n_n602_ | new_n_n611_ | new_nx0_ | new_n_n558_ | new_n_n698_ | new_n_n709_ | new_n_n601_ | new_n_n612_ | new_ng1_ | new_n_n568_ | new_n_n600_ | new_n_n609_ | new_nz0_ | new_n_n578_ | new_n_n610_ | new_n_n588_ | new_n_n599_ | new_n_n702_ | new_n_n713_ | new_n_n605_ | new_n_n616_ | new_n_n710_ | new_nw0_ | new_n_n613_ | new_n_n701_ | new_n_n711_ | new_n_n604_ | new_n_n614_ | new_n_n700_ | new_n_n699_ | new_n_n708_ | new_ny0_ | new_n_n603_;
  assign new_nd2_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_nw_ & new_n_n31_;
  assign new_n_n30_ = ~new_ny_;
  assign new_n_n23_ = ~new_nm_;
  assign new_n_n12_ = ~new_nf_;
  assign new_n_n896_ = new_n_n24_ & new_nk0_ & new_n_n30_ & new_n_n18_ & new_n_n29_ & new_n_n25_ & new_n_n21_ & new_n_n26_ & new_n_n23_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n15_;
  assign new_n_n887_ = new_n_n34_ & new_n_n10_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n20_ & new_n_n27_ & new_n_n23_ & new_n_n29_ & new_n_n30_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n797_ = new_n_n34_ & new_n_n4_ & new_n_n32_ & new_n_n33_ & new_n_n3_ & new_n_n28_ & new_n_n31_ & new_nk0_ & new_n_n15_ & new_n_n20_ & new_n_n27_ & new_n_n29_ & new_n_n30_ & new_n_n24_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n6_;
  assign new_ne2_ = new_n_n28_ & new_n_n30_ & new_nd0_ & new_n_n27_ & new_ni0_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_nw_ & new_n_n31_;
  assign new_n_n31_ = ~new_nx_;
  assign new_n_n22_ = ~new_ni0_;
  assign new_n_n13_ = ~new_ne_;
  assign new_n_n1020_ = new_n_n30_ & new_n_n27_ & new_no_ & new_n_n29_ & new_nh0_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n1009_ = new_nd0_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_n_n18_ & new_nu_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n998_ = new_nv_ & new_ni0_ & new_no_ & new_n_n30_ & new_n_n23_ & new_nh0_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n917_ = new_n_n28_ & new_n_n31_ & new_n_n22_ & new_n_n27_ & new_nj0_ & new_nk_ & new_nv_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_;
  assign new_n_n906_ = new_n_n27_ & new_n_n28_ & new_n_n15_ & new_n_n20_ & new_nk0_ & new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n25_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n807_ = new_n_n6_ & new_n_n10_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n3_ & new_n_n32_ & new_n_n20_ & new_n_n27_ & new_n_n28_ & new_n_n31_ & new_n_n30_ & new_nk0_ & new_ni0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_nb1_ = new_n_n31_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_nu_ & new_n_n18_;
  assign new_nm1_ = new_nh0_ & new_n_n24_ & new_nj0_ & new_n_n22_ & new_nz_ & new_n_n20_ & new_n_n27_ & new_n_n26_ & new_n_n25_;
  assign new_nx1_ = new_n_n28_ & new_n_n30_ & new_nd0_ & new_n_n27_ & new_ni0_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_nw_ & new_n_n31_;
  assign new_ni2_ = new_n_n25_ & new_n_n26_ & new_ni0_ & new_n_n24_ & new_nw_ & new_n_n30_ & new_n_n31_ & new_n_n27_ & new_nd0_;
  assign new_n_n25_ = ~new_nf0_;
  assign new_n_n14_ = ~new_nh0_;
  assign new_nn0_ = new_n_n916_ | new_nc1_ | new_n_n898_ | new_n_n907_ | new_n_n880_ | new_n_n889_ | new_n_n846_ | new_n_n871_ | new_n_n828_ | new_n_n837_ | new_n_n810_ | new_n_n819_ | new_n_n792_ | new_n_n801_ | new_nb1_ | new_n_n906_ | new_n_n917_ | new_n_n888_ | new_n_n899_ | new_n_n870_ | new_n_n881_ | new_n_n838_ | new_n_n856_ | new_n_n820_ | new_n_n827_ | new_n_n802_ | new_n_n809_ | new_ne1_ | new_n_n791_ | new_n_n927_ | new_n_n936_ | new_n_n900_ | new_n_n878_ | new_n_n891_ | new_n_n839_ | new_n_n869_ | new_n_n817_ | new_n_n830_ | new_n_n803_ | new_n_n808_ | new_nd1_ | new_n_n794_ | new_n_n926_ | new_n_n937_ | new_n_n890_ | new_n_n901_ | new_n_n868_ | new_n_n879_ | new_n_n840_ | new_n_n818_ | new_n_n829_ | new_n_n804_ | new_n_n807_ | new_n_n938_ | new_n_n793_ | new_n_n920_ | new_n_n929_ | new_n_n911_ | new_n_n867_ | new_n_n876_ | new_n_n832_ | new_n_n841_ | new_n_n814_ | new_n_n823_ | new_n_n788_ | new_n_n797_ | new_nf1_ | new_n_n928_ | new_n_n939_ | new_n_n910_ | new_n_n921_ | new_n_n866_ | new_n_n877_ | new_n_n813_ | new_n_n824_ | new_n_n831_ | new_n_n842_ | new_n_n940_ | new_n_n798_ | new_n_n918_ | new_n_n931_ | new_n_n896_ | new_n_n909_ | new_n_n887_ | new_n_n834_ | new_n_n843_ | new_n_n812_ | new_n_n821_ | new_n_n790_ | new_n_n799_ | new_n_n930_ | new_n_n941_ | new_n_n919_ | new_n_n897_ | new_n_n908_ | new_n_n844_ | new_n_n886_ | new_n_n822_ | new_n_n833_ | new_n_n800_ | new_n_n811_ | new_n_n789_ | new_n_n997_ | new_n_n1006_ | new_n_n979_ | new_n_n988_ | new_n_n942_ | new_n_n970_ | new_n_n924_ | new_n_n933_ | new_n_n845_ | new_n_n915_ | new_n_n996_ | new_n_n1007_ | new_n_n978_ | new_n_n989_ | new_n_n943_ | new_n_n971_ | new_n_n932_ | new_n_n914_ | new_n_n925_ | new_n_n1008_ | new_n_n835_ | new_n_n986_ | new_n_n999_ | new_n_n972_ | new_n_n977_ | new_n_n944_ | new_n_n922_ | new_n_n935_ | new_n_n825_ | new_n_n913_ | new_n_n998_ | new_n_n1009_ | new_n_n976_ | new_n_n987_ | new_n_n973_ | new_n_n934_ | new_n_n945_ | new_n_n912_ | new_n_n923_ | new_nh1_ | new_n_n815_ | new_n_n1010_ | new_nt1_ | new_n_n992_ | new_n_n1001_ | new_n_n966_ | new_n_n983_ | new_n_n893_ | new_n_n902_ | new_n_n875_ | new_n_n884_ | new_n_n805_ | new_nv1_ | new_ng1_ | new_n_n1000_ | new_n_n1011_ | new_n_n982_ | new_n_n993_ | new_n_n903_ | new_n_n967_ | new_n_n885_ | new_n_n892_ | new_n_n795_ | new_n_n874_ | new_n_n1025_ | new_nf2_ | new_n_n1003_ | new_n_n1012_ | new_n_n990_ | new_n_n968_ | new_n_n981_ | new_n_n1024_ | new_ne2_ | new_n_n1002_ | new_n_n1013_ | new_n_n873_ | new_n_n882_ | new_n_n895_ | new_n_n904_ | new_n_n980_ | new_n_n991_ | new_n_n905_ | new_n_n969_ | new_n_n883_ | new_n_n894_ | new_n_n872_ | new_ny1_ | new_nl1_ | new_n_n1005_ | new_n_n1014_ | new_n_n1023_ | new_nh2_ | new_nz1_ | new_nk1_ | new_ng2_ | new_n_n1015_ | new_n_n1022_ | new_nj1_ | new_n_n1004_ | new_nj2_ | new_nw1_ | new_n_n994_ | new_n_n1021_ | new_n_n985_ | new_nx1_ | new_ni1_ | new_nc2_ | new_ns1_ | new_n_n1019_ | new_n_n1028_ | new_n_n984_ | new_n_n995_ | new_n_n1020_ | new_ni2_ | new_n_n964_ | new_n_n974_ | new_nq1_ | new_n_n955_ | new_n_n1029_ | new_nd2_ | new_n_n1018_ | new_n_n965_ | new_n_n975_ | new_np1_ | new_n_n954_ | new_n_n1026_ | new_na2_ | new_n_n962_ | new_n_n1017_ | new_n_n953_ | new_nm1_ | new_n_n865_ | new_n_n1027_ | new_nb2_ | new_n_n963_ | new_n_n1016_ | new_n_n855_ | new_n_n952_ | new_n_n960_ | new_n_n863_ | new_n_n951_ | new_n_n961_ | new_n_n854_ | new_n_n864_ | new_n_n950_ | new_nw0_ | new_n_n853_ | new_n_n949_ | new_n_n958_ | new_n_n852_ | new_n_n861_ | new_n_n948_ | new_n_n959_ | new_n_n851_ | new_n_n862_ | new_n_n796_ | new_n_n956_ | new_ny0_ | new_na1_ | new_n_n816_ | new_n_n848_ | new_n_n857_ | new_nz0_ | new_n_n826_ | new_n_n858_ | new_n_n836_ | new_n_n847_ | new_n_n859_ | new_n_n947_ | new_n_n806_ | new_n_n850_ | new_n_n957_ | new_nx0_ | new_n_n946_ | new_n_n849_ | new_n_n860_;
  assign new_n_n1021_ = new_n_n29_ & new_n_n30_ & new_n_n26_ & new_n_n25_ & new_nu_ & new_n_n27_ & new_n_n22_ & new_nd0_ & new_n_n24_ & new_n_n18_;
  assign new_n_n1008_ = new_nd0_ & new_n_n27_ & new_n_n18_ & new_ni0_ & new_n_n30_ & new_nu_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n999_ = new_nj0_ & new_n_n22_ & new_no_ & new_nv_ & new_n_n23_ & new_nh0_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n916_ = new_n_n22_ & new_n_n27_ & new_nd_ & new_nj0_ & new_n_n5_ & new_nk_ & new_nv_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n31_ & new_n_n28_;
  assign new_n_n907_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_n_n15_ & new_n_n30_ & new_nk0_ & new_n_n26_ & new_n_n25_ & new_n_n10_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n817_ = new_n_n32_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_ni0_ & new_n_n20_ & new_n_n21_ & new_n_n30_ & new_nk0_ & new_n_n15_ & new_n_n25_ & new_n_n7_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_nc1_ = new_n_n31_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n23_ & new_n_n33_ & new_n_n34_ & new_nu_ & new_n_n18_;
  assign new_nl1_ = new_n_n28_ & new_nz_ & new_n_n20_ & new_n_n27_ & new_nh0_ & new_ni0_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_ny1_ = new_n_n29_ & new_nz_ & new_n_n27_ & new_n_n28_ & new_nh0_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_n_n31_ & new_n_n30_;
  assign new_nh2_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_n_n23_ & new_n_n33_ & new_n_n34_ & new_nw_ & new_n_n31_;
  assign new_n_n24_ = ~new_ng0_;
  assign new_n_n15_ = ~new_nj0_;
  assign new_n_n1029_ = new_n_n24_ & new_nk0_ & new_n_n26_ & new_n_n25_ & new_n_n1_ & new_n_n20_ & new_n_n27_ & new_n_n22_ & new_nj0_;
  assign new_n_n1018_ = new_no_ & new_n_n30_ & new_n_n26_ & new_n_n25_ & new_nh0_ & new_n_n31_ & new_ni0_ & new_n_n27_ & new_n_n24_ & new_nv_;
  assign new_n_n1011_ = new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_nf0_ & new_n_n23_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n31_;
  assign new_n_n1000_ = new_ni0_ & new_n_n27_ & new_n_n30_ & new_nv_ & new_no_ & new_nh0_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n937_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_nk0_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n31_ & new_n_n28_;
  assign new_n_n926_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n20_ & new_nj0_ & new_n_n5_ & new_nd_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n827_ = new_n_n34_ & new_n_n6_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_n_n18_ & new_nk0_ & new_nd0_ & new_n_n2_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n10_;
  assign new_n_n49_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n9_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n38_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_nz1_ = new_n_n25_ & new_n_n26_ & new_nh0_ & new_n_n24_ & new_ni0_ & new_no_ & new_n_n30_ & new_n_n31_ & new_n_n27_ & new_n_n20_;
  assign new_n_n34_ = ~new_nn_;
  assign new_n_n27_ = ~new_nc0_;
  assign new_n_n16_ = ~new_nc_;
  assign new_n_n1028_ = new_n_n25_ & new_n_n18_ & new_nu_ & new_n_n26_ & new_n_n27_ & new_n_n22_ & new_nd0_ & new_nj0_ & new_n_n24_;
  assign new_n_n1019_ = new_n_n29_ & new_n_n30_ & new_n_n23_ & new_no_ & new_nh0_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n1010_ = new_n_n30_ & new_n_n27_ & new_n_n21_ & new_n_n29_ & new_nf0_ & new_n_n23_ & new_nh_ & new_n_n33_ & new_n_n6_ & new_n_n31_ & new_n_n28_;
  assign new_n_n1001_ = new_n_n22_ & new_n_n27_ & new_nv_ & new_nj0_ & new_no_ & new_nh0_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n936_ = new_n_n22_ & new_n_n20_ & new_nk0_ & new_nj0_ & new_n_n24_ & new_n_n23_ & new_n_n21_ & new_n_n26_ & new_n_n1_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n927_ = new_n_n31_ & new_n_n3_ & new_n_n27_ & new_n_n28_ & new_n_n20_ & new_nj0_ & new_n_n22_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n32_;
  assign new_n_n837_ = new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n32_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n30_ & new_n_n18_ & new_n_n24_ & new_nk0_ & new_n_n21_ & new_n_n29_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n1_ & new_n_n6_;
  assign new_n_n48_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n39_ = new_n_n15_ & new_n_n27_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_na2_ = new_n_n29_ & new_nz_ & new_n_n27_ & new_n_n28_ & new_nh0_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n30_;
  assign new_nj2_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_nw_ & new_n_n31_;
  assign new_n_n26_ = ~new_ne0_;
  assign new_n_n17_ = ~new_nu_;
  assign new_n_n991_ = new_n_n18_ & new_nd0_ & new_n_n29_ & new_n_n30_ & new_n_n23_ & new_na_ & new_n_n34_ & new_n_n31_ & new_n_n33_ & new_n_n28_ & new_n_n27_;
  assign new_n_n980_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n20_ & new_nj0_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n31_;
  assign new_n_n969_ = new_n_n31_ & new_n_n3_ & new_n_n27_ & new_n_n28_ & new_n_n30_ & new_nk_ & new_n_n29_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n4_ & new_n_n33_ & new_n_n32_;
  assign new_n_n958_ = new_ni0_ & new_n_n27_ & new_n_n30_ & new_nv_ & new_n_n21_ & new_nf0_ & new_nk_ & new_n_n23_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n28_;
  assign new_n_n957_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_n_n22_ & new_nk0_ & new_nj0_ & new_n_n26_ & new_n_n1_ & new_n_n34_ & new_n_n10_ & new_n_n33_ & new_n_n32_;
  assign new_n_n946_ = new_n_n20_ & new_n_n27_ & new_n_n24_ & new_nk0_ & new_n_n30_ & new_n_n21_ & new_n_n29_ & new_n_n26_ & new_n_n1_ & new_n_n32_ & new_n_n33_ & new_n_n31_ & new_n_n28_;
  assign new_n_n847_ = new_n_n6_ & new_n_n10_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n28_ & new_n_n31_ & new_nj0_ & new_n_n22_ & new_n_n20_ & new_n_n27_ & new_n_n21_ & new_nk0_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n1_;
  assign new_n_n50_ = new_n_n29_ & new_n_n8_ & new_n_n24_ & new_n_n27_ & new_n_n15_ & new_n_n13_ & new_nm0_ & new_n_n9_ & new_n_n20_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n47_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_n_n20_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_nl_ & new_nj_ & new_n_n34_ & new_n_n30_;
  assign new_n_n36_ = new_n_n15_ & new_n_n27_ & new_n_n13_ & new_nm0_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_nf1_ = new_n_n27_ & new_n_n28_ & new_nh0_ & new_n_n20_ & new_n_n22_ & new_nj0_ & new_n_n34_ & new_n_n33_ & new_no_ & new_n_n32_ & new_n_n31_;
  assign new_nq1_ = new_n_n25_ & new_n_n26_ & new_nh0_ & new_n_n24_ & new_ni0_ & new_n_n31_ & new_nz_ & new_n_n30_ & new_n_n27_ & new_n_n20_;
  assign new_n_n29_ = ~new_na0_;
  assign new_n_n18_ = ~new_nv_;
  assign new_n_n990_ = new_n_n30_ & new_n_n18_ & new_n_n21_ & new_n_n29_ & new_n_n23_ & new_na_ & new_n_n33_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_nd0_;
  assign new_n_n981_ = new_n_n27_ & new_n_n28_ & new_n_n29_ & new_n_n30_ & new_n_n21_ & new_nf0_ & new_nk_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n32_ & new_n_n31_;
  assign new_n_n968_ = new_n_n27_ & new_n_n28_ & new_n_n5_ & new_nd_ & new_n_n30_ & new_nk_ & new_n_n29_ & new_nf0_ & new_nh_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n959_ = new_n_n20_ & new_n_n27_ & new_n_n30_ & new_ni0_ & new_n_n21_ & new_nf0_ & new_nk_ & new_n_n23_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n28_;
  assign new_n_n956_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_n_n20_ & new_nj0_ & new_n_n24_ & new_nk0_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n34_ & new_n_n32_ & new_n_n31_;
  assign new_n_n947_ = new_n_n27_ & new_n_n28_ & new_nk0_ & new_n_n20_ & new_n_n30_ & new_n_n21_ & new_n_n29_ & new_n_n26_ & new_n_n1_ & new_n_n33_ & new_n_n10_ & new_n_n32_ & new_n_n31_;
  assign new_n_n857_ = new_n_n33_ & new_n_n34_ & new_n_n28_ & new_n_n31_ & new_n_n27_ & new_n_n15_ & new_n_n20_ & new_n_n25_ & new_n_n29_ & new_n_n30_ & new_nk0_ & new_n_n23_ & new_n_n16_ & new_n_n12_ & new_n_n13_ & new_n_n11_ & new_n_n10_;
  assign new_n_n51_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n46_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n37_ = new_n_n15_ & new_n_n24_ & new_n_n14_ & new_nm0_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n27_;
  assign new_ng1_ = new_n_n27_ & new_n_n28_ & new_n_n22_ & new_nd0_ & new_nj0_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_nw_ & new_n_n31_;
  assign new_np1_ = new_n_n25_ & new_n_n26_ & new_nh0_ & new_n_n24_ & new_n_n22_ & new_n_n30_ & new_n_n29_ & new_nz_ & new_n_n27_ & new_n_n20_;
  assign new_n_n28_ = ~new_nb0_;
  assign new_n_n19_ = ~new_nw_;
  assign new_n_n989_ = new_n_n28_ & new_n_n31_ & new_n_n20_ & new_n_n27_ & new_n_n22_ & new_nf0_ & new_nj0_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n978_ = new_n_n27_ & new_n_n28_ & new_ni0_ & new_n_n20_ & new_n_n30_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n31_;
  assign new_n_n971_ = new_n_n28_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n21_ & new_nc_ & new_nn_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n960_ = new_n_n22_ & new_n_n27_ & new_nv_ & new_nj0_ & new_n_n21_ & new_nf0_ & new_nk_ & new_n_n23_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n28_;
  assign new_n_n52_ = new_n_n29_ & new_n_n8_ & new_n_n15_ & new_n_n27_ & new_nm0_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_nt_ & new_n_n10_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n45_ = new_n_n24_ & new_n_n27_ & new_nm0_ & new_n_n15_ & new_n_n14_ & new_n_n12_ & new_n_n13_ & new_n_n9_ & new_n_n20_ & new_nt_ & new_n_n11_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n29_;
  assign new_nw0_ = new_n_n31_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_nc_ & new_n_n21_ & new_n_n23_ & new_n_n33_ & new_n_n17_;
  assign new_nd1_ = new_n_n31_ & new_n_n19_ & new_n_n29_ & new_n_n30_ & new_n_n28_ & new_nd0_ & new_n_n27_ & new_n_n34_ & new_n_n32_ & new_n_n33_ & new_nu_ & new_n_n18_;
  assign new_no1_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nd0_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_nv_ & new_n_n19_;
  assign new_nv1_ = new_n_n28_ & new_n_n30_ & new_n_n20_ & new_n_n27_ & new_nh0_ & new_ni0_ & new_n_n34_ & new_n_n33_ & new_no_ & new_n_n32_ & new_n_n31_;
  assign new_ng2_ = new_n_n25_ & new_n_n26_ & new_n_n22_ & new_n_n24_ & new_nw_ & new_n_n29_ & new_n_n30_ & new_n_n27_ & new_nd0_;
  assign new_n_n988_ = new_n_n28_ & new_n_n31_ & new_n_n22_ & new_n_n27_ & new_nj0_ & new_nf0_ & new_nv_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n979_ = new_n_n27_ & new_n_n28_ & new_nj0_ & new_n_n22_ & new_nv_ & new_n_n23_ & new_nf0_ & new_nh_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n31_;
  assign new_n_n970_ = new_n_n28_ & new_n_n31_ & new_nd0_ & new_n_n27_ & new_n_n18_ & new_n_n29_ & new_n_n30_ & new_n_n2_ & new_nc_ & new_n_n34_ & new_n_n6_ & new_n_n33_ & new_n_n32_;
  assign new_n_n961_ = new_n_n20_ & new_n_n27_ & new_nj0_ & new_n_n22_ & new_n_n21_ & new_nf0_ & new_nk_ & new_n_n23_ & new_nh_ & new_n_n33_ & new_nn_ & new_n_n31_ & new_n_n28_;
  assign new_n_n53_ = new_n_n27_ & new_n_n29_ & new_n_n15_ & new_n_n24_ & new_nm0_ & new_n_n13_ & new_n_n14_ & new_n_n9_ & new_nt_ & new_n_n11_ & new_n_n12_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n19_ & new_n_n30_;
  assign new_n_n44_ = new_n_n27_ & new_n_n29_ & new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n11_ & new_n_n12_ & new_n_n9_ & new_n_n20_ & new_nt_ & new_n_n10_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n8_;
  assign new_n_n35_ = new_nm0_ & new_n_n15_ & new_n_n13_ & new_n_n14_ & new_n_n12_ & new_n_n10_ & new_n_n11_ & new_n_n9_ & new_ni0_ & new_n_n20_ & new_nt_ & new_n_n23_ & new_n_n16_ & new_n_n34_ & new_nj_ & new_n_n30_ & new_n_n27_;
  assign new_ne1_ = new_n_n27_ & new_n_n28_ & new_nh0_ & new_n_n20_ & new_n_n22_ & new_nj0_ & new_n_n23_ & new_no_ & new_n_n34_ & new_n_n33_ & new_n_n31_;
  assign new_nn1_ = new_n_n30_ & new_n_n31_ & new_n_n28_ & new_n_n29_ & new_n_n27_ & new_nd0_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_nv_ & new_n_n19_;
  assign new_nw1_ = new_n_n28_ & new_n_n30_ & new_nd0_ & new_n_n27_ & new_ni0_ & new_n_n23_ & new_n_n33_ & new_n_n21_ & new_nw_ & new_n_n31_;
  assign new_nf2_ = new_n_n29_ & new_n_n30_ & new_n_n27_ & new_n_n28_ & new_nd0_ & new_n_n21_ & new_n_n32_ & new_n_n33_ & new_nw_ & new_n_n31_;
endmodule


