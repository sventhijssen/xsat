// Benchmark "top" written by ABC on Fri Mar 31 12:11:20 2023

module top ( 
    txwrd3, a, qpr4, txwrd2, b, i1zzz0, txwrd5, c, p1zzz0, txwrd4, xzfs,
    i1zzz2, i2zzz1, p1zzz1, p2zzz0, qpr1, i1zzz1, i2zzz0, p1zzz2, p2zzz1,
    qpr0, i1zzz4, i2zzz3, infin, p1zzz3, p2zzz2, qpr3, txwrd1, vybb1,
    i1zzz3, i2zzz2, p1zzz4, p2zzz3, qpr2, txwrd0, vybb0, comppar, psrw,
    xz323, cbt2, mmerr, ryz, xz324, esrsum, v1zzz7, v2zzz6, xz161, pfin,
    stw_n, v2zzz7, vzzze, xz162, xz320, cbt1, slad0, v1zzz5, v2zzz4, xz163,
    xz321, cbt0, slad1, v1zzz6, v2zzz5, xz322, pybb5, slad2, txwrd14,
    v1zzz3, v2zzz2, xz160_n, pybb4, slad3, txwrd13, v1zzz4, v2zzz3, iclr,
    pybb3, rptwin, txwrd12, v1zzz1, v2zzz0, pybb2, txwrd11, v1zzz2, v2zzz1,
    axz1, inzzze, axz0, pybb8, v1zzz0, inybb8, pybb7, xzfr0, enwin, ofs1,
    pybb6, pzzze, txmess_n, txwrd15, xzfr1, i1zzz6, i2zzz5, inybb6, ofs2,
    p1zzz5, p2zzz4, rxz0, i1zzz5, i2zzz4, inybb7, p1zzz6, p2zzz5, rpten,
    rxz1, i2zzz7, inybb4, p1zzz7, p2zzz6, i1zzz7, i2zzz6, inybb5, p2zzz7,
    inybb2, pybb1, txwrd7, txwrd10, inybb3, pybb0, txwrd6, inybb0, txwrd9,
    inybb1, psync, txwrd8, vfin,
    i1zzz0_p, v1zzz0_p, i1zzz3_p, i2zzz2_p, txwrd8_p, v1zzz2_p, v2zzz1_p,
    i1zzz4_p, i2zzz3_p, stw_f, txwrd9_p, v1zzz1_p, v2zzz0_p, xz163_p, c_p,
    enwin_p, i1zzz1_p, i2zzz0_p, txwrd6_p, v1zzz4_p, v2zzz3_p, i1zzz2_p,
    i2zzz1_p, txwrd7_p, v1zzz3_p, v2zzz2_p, p1zzz4_p, p2zzz3_p, xz162_p,
    b_p, p1zzz3_p, p2zzz2_p, p1zzz2_p, p2zzz1_p, xzfr1_p, p1zzz1_p,
    p2zzz0_p, txwrd14_p, xz161_p, a_p, p1zzz0_p, axz0_p, txwrd15_p, axz1_p,
    td_p, fsesr_p, rptwin_p, txwrd12_p, txwrd11_p, xz322_p, p2zzz7_p,
    txwrd13_p, xz324_p, xzfs_p, p1zzz7_p, p2zzz6_p, xzfr0_p, p1zzz6_p,
    p2zzz5_p, rxz1_p, comppar_p, ofs2_p, p1zzz5_p, p2zzz4_p, rxz0_p,
    xz323_p, i1zzz7_p, i2zzz6_p, ofs1_p, ryz_p, sbuff, txwrd4_p, v1zzz6_p,
    v2zzz5_p, xz160_f, xz320_p, i2zzz7_p, txwrd5_p, v1zzz5_p, v2zzz4_p,
    i1zzz5_p, i2zzz4_p, qpr4_p, txwrd2_p, v2zzz7_p, i1zzz6_p, i2zzz5_p,
    txwrd3_p, v1zzz7_p, v2zzz6_p, qpr2_p, txwrd0_p, qpr3_p, txwrd1_p,
    xz321_p, qpr0_p, qpr1_p, txmess_f, txwrd10_p  );
  input  txwrd3, a, qpr4, txwrd2, b, i1zzz0, txwrd5, c, p1zzz0, txwrd4,
    xzfs, i1zzz2, i2zzz1, p1zzz1, p2zzz0, qpr1, i1zzz1, i2zzz0, p1zzz2,
    p2zzz1, qpr0, i1zzz4, i2zzz3, infin, p1zzz3, p2zzz2, qpr3, txwrd1,
    vybb1, i1zzz3, i2zzz2, p1zzz4, p2zzz3, qpr2, txwrd0, vybb0, comppar,
    psrw, xz323, cbt2, mmerr, ryz, xz324, esrsum, v1zzz7, v2zzz6, xz161,
    pfin, stw_n, v2zzz7, vzzze, xz162, xz320, cbt1, slad0, v1zzz5, v2zzz4,
    xz163, xz321, cbt0, slad1, v1zzz6, v2zzz5, xz322, pybb5, slad2,
    txwrd14, v1zzz3, v2zzz2, xz160_n, pybb4, slad3, txwrd13, v1zzz4,
    v2zzz3, iclr, pybb3, rptwin, txwrd12, v1zzz1, v2zzz0, pybb2, txwrd11,
    v1zzz2, v2zzz1, axz1, inzzze, axz0, pybb8, v1zzz0, inybb8, pybb7,
    xzfr0, enwin, ofs1, pybb6, pzzze, txmess_n, txwrd15, xzfr1, i1zzz6,
    i2zzz5, inybb6, ofs2, p1zzz5, p2zzz4, rxz0, i1zzz5, i2zzz4, inybb7,
    p1zzz6, p2zzz5, rpten, rxz1, i2zzz7, inybb4, p1zzz7, p2zzz6, i1zzz7,
    i2zzz6, inybb5, p2zzz7, inybb2, pybb1, txwrd7, txwrd10, inybb3, pybb0,
    txwrd6, inybb0, txwrd9, inybb1, psync, txwrd8, vfin;
  output i1zzz0_p, v1zzz0_p, i1zzz3_p, i2zzz2_p, txwrd8_p, v1zzz2_p, v2zzz1_p,
    i1zzz4_p, i2zzz3_p, stw_f, txwrd9_p, v1zzz1_p, v2zzz0_p, xz163_p, c_p,
    enwin_p, i1zzz1_p, i2zzz0_p, txwrd6_p, v1zzz4_p, v2zzz3_p, i1zzz2_p,
    i2zzz1_p, txwrd7_p, v1zzz3_p, v2zzz2_p, p1zzz4_p, p2zzz3_p, xz162_p,
    b_p, p1zzz3_p, p2zzz2_p, p1zzz2_p, p2zzz1_p, xzfr1_p, p1zzz1_p,
    p2zzz0_p, txwrd14_p, xz161_p, a_p, p1zzz0_p, axz0_p, txwrd15_p, axz1_p,
    td_p, fsesr_p, rptwin_p, txwrd12_p, txwrd11_p, xz322_p, p2zzz7_p,
    txwrd13_p, xz324_p, xzfs_p, p1zzz7_p, p2zzz6_p, xzfr0_p, p1zzz6_p,
    p2zzz5_p, rxz1_p, comppar_p, ofs2_p, p1zzz5_p, p2zzz4_p, rxz0_p,
    xz323_p, i1zzz7_p, i2zzz6_p, ofs1_p, ryz_p, sbuff, txwrd4_p, v1zzz6_p,
    v2zzz5_p, xz160_f, xz320_p, i2zzz7_p, txwrd5_p, v1zzz5_p, v2zzz4_p,
    i1zzz5_p, i2zzz4_p, qpr4_p, txwrd2_p, v2zzz7_p, i1zzz6_p, i2zzz5_p,
    txwrd3_p, v1zzz7_p, v2zzz6_p, qpr2_p, txwrd0_p, qpr3_p, txwrd1_p,
    xz321_p, qpr0_p, qpr1_p, txmess_f, txwrd10_p;
  wire new_ntxwrd3_, new_na_, new_nqpr4_, new_ntxwrd2_, new_nb_,
    new_ni1zzz0_, new_ntxwrd5_, new_nc_, new_np1zzz0_, new_ntxwrd4_,
    new_nxzfs_, new_ni1zzz2_, new_ni2zzz1_, new_np1zzz1_, new_np2zzz0_,
    new_nqpr1_, new_ni1zzz1_, new_ni2zzz0_, new_np1zzz2_, new_np2zzz1_,
    new_nqpr0_, new_ni1zzz4_, new_ni2zzz3_, new_ninfin_, new_np1zzz3_,
    new_np2zzz2_, new_nqpr3_, new_ntxwrd1_, new_nvybb1_, new_ni1zzz3_,
    new_ni2zzz2_, new_np1zzz4_, new_np2zzz3_, new_nqpr2_, new_ntxwrd0_,
    new_nvybb0_, new_ncomppar_, new_npsrw_, new_nxz323_, new_ncbt2_,
    new_nmmerr_, new_nryz_, new_nxz324_, new_nesrsum_, new_nv1zzz7_,
    new_nv2zzz6_, new_nxz161_, new_npfin_, new_nstw_n_, new_nv2zzz7_,
    new_nvzzze_, new_nxz162_, new_nxz320_, new_ncbt1_, new_nslad0_,
    new_nv1zzz5_, new_nv2zzz4_, new_nxz163_, new_nxz321_, new_ncbt0_,
    new_nslad1_, new_nv1zzz6_, new_nv2zzz5_, new_nxz322_, new_npybb5_,
    new_nslad2_, new_ntxwrd14_, new_nv1zzz3_, new_nv2zzz2_, new_nxz160_n_,
    new_npybb4_, new_nslad3_, new_ntxwrd13_, new_nv1zzz4_, new_nv2zzz3_,
    new_niclr_, new_npybb3_, new_nrptwin_, new_ntxwrd12_, new_nv1zzz1_,
    new_nv2zzz0_, new_npybb2_, new_ntxwrd11_, new_nv1zzz2_, new_nv2zzz1_,
    new_naxz1_, new_ninzzze_, new_naxz0_, new_npybb8_, new_nv1zzz0_,
    new_ninybb8_, new_npybb7_, new_nxzfr0_, new_nenwin_, new_nofs1_,
    new_npybb6_, new_npzzze_, new_ntxmess_n_, new_ntxwrd15_, new_nxzfr1_,
    new_ni1zzz6_, new_ni2zzz5_, new_ninybb6_, new_nofs2_, new_np1zzz5_,
    new_np2zzz4_, new_nrxz0_, new_ni1zzz5_, new_ni2zzz4_, new_ninybb7_,
    new_np1zzz6_, new_np2zzz5_, new_nrpten_, new_nrxz1_, new_ni2zzz7_,
    new_ninybb4_, new_np1zzz7_, new_np2zzz6_, new_ni1zzz7_, new_ni2zzz6_,
    new_ninybb5_, new_np2zzz7_, new_ninybb2_, new_npybb1_, new_ntxwrd7_,
    new_ntxwrd10_, new_ninybb3_, new_npybb0_, new_ntxwrd6_, new_ninybb0_,
    new_ntxwrd9_, new_ninybb1_, new_npsync_, new_ntxwrd8_, new_nvfin_,
    new_nsbuff_, new_n_n378_, new_np1zzz5_p_, new_n_n363_, new_n_n356_,
    new_ni1zzz0_p_, new_n_n341_, new_n_n334_, new_ni2zzz3_p_, new_n_n319_,
    new_nxzfr1_p_, new_nofs1_p_, new_n_n304_, new_n_n298_, new_nv1zzz4_p_,
    new_n_n283_, new_n_n276_, new_nv2zzz7_p_, new_n_n262_, new_ntxwrd6_p_,
    new_n_n246_, new_nxz323_p_, new_n_n226_, new_nmis16706_,
    new_nmis11584_, new_n_n212_, new_nmis16544_, new_n_n201_, new_n_n197_,
    new_n_n178_, new_nmis16631_, new_n_n161_, new_n_n153_, new_nmis11560_,
    new_nmis10125_, new_nmis16690_, new_nmis9174_, new_n_n109_,
    new_n_n105_, new_nmis16742_, new_nmis9255_, new_nmis16866_,
    new_n_n371_, new_n_n370_, new_n_n364_, new_n_n355_, new_n_n349_,
    new_ni1zzz4_p_, new_ni1zzz7_p_, new_n_n326_, new_n_n320_, new_n_n314_,
    new_nofs2_p_, new_na_p_, new_n_n297_, new_n_n291_, new_nv2zzz0_p_,
    new_nv2zzz3_p_, new_n_n268_, new_ntxwrd3_p_, new_n_n253_, new_n_n247_,
    new_n_n233_, new_n_n227_, new_n_n220_, new_nmis11583_, new_nmis8027_,
    new_n_n208_, new_n_n200_, new_nmis16553_, new_nmis16726_, new_n_n169_,
    new_n_n162_, new_n_n152_, new_n_n145_, new_nmis9071_, new_n_n136_,
    new_n_n113_, new_n_n110_, new_n_n104_, new_n_n97_, new_nmis16577_,
    new_n_n85_, new_n_n379_, new_n_n372_, new_np2zzz5_p_, new_n_n347_,
    new_ni1zzz3_p_, new_n_n335_, new_n_n325_, new_n_n318_, new_n_n316_,
    new_n_n309_, new_nv1zzz1_p_, new_n_n289_, new_nv1zzz7_p_, new_n_n277_,
    new_n_n267_, new_n_n260_, new_n_n255_, new_ntxwrd9_p_, new_n_n232_,
    new_n_n225_, new_nmis16790_, new_nmis11582_, new_nmis15083_,
    new_nmis16541_, new_n_n202_, new_n_n198_, new_n_n184_, new_n_n176_,
    new_nmis16609_, new_n_n151_, new_n_n144_, new_nmis16754_, new_n_n137_,
    new_n_n123_, new_n_n118_, new_n_n103_, new_nmis16778_, new_n_n92_,
    new_n_n86_, new_nstw_f_, new_np1zzz1_p_, new_np1zzz4_p_, new_n_n354_,
    new_n_n348_, new_n_n342_, new_n_n336_, new_ni2zzz4_p_, new_ni2zzz7_p_,
    new_n_n315_, new_n_n310_, new_n_n296_, new_n_n290_, new_n_n284_,
    new_n_n278_, new_ntxwrd0_p_, new_n_n261_, new_n_n254_, new_n_n248_,
    new_nxz324_p_, new_nxz162_p_, new_n_n221_, new_nmis11581_,
    new_nmis16613_, new_n_n207_, new_nmis16762_, new_n_n199_, new_n_n183_,
    new_n_n177_, new_n_n170_, new_nmis16736_, new_nmis15339_, new_n_n141_,
    new_nmis16786_, new_nmis16724_, new_n_n119_, new_nmis16598_,
    new_nmis16604_, new_n_n91_, new_nmis16864_, new_n_n368_,
    new_np2zzz2_p_, new_n_n344_, new_ni1zzz6_p_, new_nqpr0_p_, new_n_n301_,
    new_nv2zzz2_p_, new_ntxwrd1_p_, new_ntxwrd13_p_, new_nxz320_p_,
    new_n_n211_, new_n_n205_, new_nmis11591_, new_n_n190_, new_n_n150_,
    new_nmis16730_, new_nmis16588_, new_n_n133_, new_nmis11154_,
    new_n_n102_, new_n_n95_, new_nmis16579_, new_nmis16670_, new_n_n9_,
    new_n_n367_, new_n_n361_, new_n_n343_, new_n_n337_, new_n_n308_,
    new_n_n302_, new_n_n285_, new_ntxwrd4_p_, new_n_n245_, new_n_n238_,
    new_nmis16879_, new_n_n206_, new_nmis11592_, new_n_n191_, new_n_n149_,
    new_nmis11578_, new_nmis16701_, new_n_n132_, new_nmis16887_,
    new_n_n101_, new_n_n96_, new_n_n88_, new_nmis16665_, new_n_n369_,
    new_n_n362_, new_n_n357_, new_n_n350_, new_nb_p_, new_nqpr3_p_,
    new_n_n292_, new_n_n252_, new_ntxwrd11_p_, new_n_n239_, new_nmis16629_,
    new_nmis11589_, new_n_n192_, new_n_n148_, new_n_n140_, new_n_n134_,
    new_n_n100_, new_n_n94_, new_n_n90_, new_n_n83_, new_np1zzz6_p_,
    new_np2zzz1_p_, new_np2zzz4_p_, new_np2zzz7_p_, new_nc_p_, new_n_n303_,
    new_nv1zzz0_p_, new_ntxwrd10_p_, new_ntxwrd12_p_, new_ntxwrd15_p_,
    new_nmis16581_, new_n_n196_, new_nmis11590_, new_n_n143_,
    new_nmis15848_, new_n_n135_, new_nmis16625_, new_nmis16780_,
    new_n_n89_, new_n_n84_, new_ntd_p_, new_n_n376_, new_n_n365_,
    new_n_n358_, new_n_n317_, new_nxzfs_p_, new_n_n306_, new_naxz0_p_,
    new_nv1zzz3_p_, new_n_n251_, new_ntxwrd14_p_, new_nxz322_p_,
    new_n_n228_, new_nmis11547_, new_n_n194_, new_n_n187_, new_n_n180_,
    new_n_n172_, new_n_n163_, new_nmis16712_, new_n_n126_, new_nmis15964_,
    new_nmis8768_, new_nmis16593_, new_n_n107_, new_n_n5_, new_nfsesr_p_,
    new_np1zzz2_p_, new_np2zzz0_p_, new_np2zzz3_p_, new_ntxmess_f_,
    new_n_n313_, new_n_n305_, new_n_n299_, new_n_n286_, new_n_n259_,
    new_n_n242_, new_n_n236_, new_nxz161_p_, new_nenwin_p_, new_n_n193_,
    new_n_n188_, new_n_n179_, new_nmis16618_, new_n_n156_, new_n_n130_,
    new_nmis16565_, new_n_n122_, new_n_n115_, new_n_n111_, new_n_n108_,
    new_n_n6_, new_n_n377_, new_np1zzz7_p_, new_n_n359_, new_ni2zzz1_p_,
    new_n_n323_, new_n_n307_, new_n_n300_, new_n_n279_, new_n_n266_,
    new_n_n244_, new_n_n237_, new_nmis11585_, new_n_n215_, new_nmis16591_,
    new_nmis16585_, new_nmis16732_, new_n_n165_, new_nmis16623_,
    new_nmis16710_, new_n_n127_, new_n_n121_, new_n_n114_, new_nmis16893_,
    new_nmis16620_, new_n_n7_, new_n_n383_, new_n_n366_, new_n_n360_,
    new_n_n330_, new_n_n324_, new_nqpr1_p_, new_nqpr4_p_, new_nv2zzz5_p_,
    new_n_n272_, new_n_n243_, new_nxz321_p_, new_nmis11586_, new_n_n216_,
    new_n_n195_, new_n_n189_, new_n_n171_, new_n_n164_, new_n_n157_,
    new_n_n131_, new_n_n128_, new_n_n120_, new_nmis16758_, new_nmis11546_,
    new_nmis11549_, new_n_n8_, new_np1zzz0_p_, new_n_n373_, new_n_n353_,
    new_n_n346_, new_ni1zzz5_p_, new_n_n331_, new_n_n329_, new_n_n322_,
    new_nrptwin_p_, new_nrxz1_p_, new_n_n295_, new_n_n288_, new_nv2zzz1_p_,
    new_n_n273_, new_n_n271_, new_ntxwrd2_p_, new_ntxwrd5_p_, new_n_n249_,
    new_n_n231_, new_nxz163_p_, new_nmis11587_, new_n_n217_,
    new_nmis16722_, new_nmis16788_, new_nmis16760_, new_nmis16615_,
    new_nmis16606_, new_n_n182_, new_n_n175_, new_nmis16627_, new_n_n158_,
    new_nmis16583_, new_nmis16740_, new_n_n138_, new_nmis16885_,
    new_nmis7401_, new_nmis15650_, new_n_n116_, new_nmis16555_,
    new_nmis11548_, new_n_n93_, new_nmis16858_, new_n_n1_, new_n_n380_,
    new_n_n374_, new_np2zzz6_p_, new_ni1zzz1_p_, new_n_n338_, new_n_n332_,
    new_ni2zzz2_p_, new_ni2zzz5_p_, new_nxzfr0_p_, new_n_n311_,
    new_nv1zzz2_p_, new_nv1zzz5_p_, new_n_n280_, new_n_n274_,
    new_nv2zzz6_p_, new_n_n265_, new_n_n256_, new_n_n250_, new_n_n230_,
    new_n_n224_, new_nmis11588_, new_nmis16569_, new_n_n214_, new_n_n210_,
    new_n_n203_, new_nmis16546_, new_nmis15081_, new_nmis15080_,
    new_nmis16633_, new_n_n166_, new_n_n159_, new_n_n155_, new_n_n142_,
    new_nmis16602_, new_nmis16891_, new_n_n124_, new_nmis15847_,
    new_n_n117_, new_nmis16889_, new_nmis11562_, new_nmis16716_,
    new_n_n87_, new_n_n2_, new_n_n382_, new_np1zzz3_p_, new_n_n352_,
    new_ni1zzz2_p_, new_n_n340_, new_ni2zzz0_p_, new_n_n328_,
    new_ni2zzz6_p_, new_nryz_p_, new_n_n312_, new_nqpr2_p_, new_n_n294_,
    new_nv1zzz6_p_, new_n_n282_, new_nv2zzz4_p_, new_n_n270_, new_n_n263_,
    new_n_n258_, new_ntxwrd8_p_, new_n_n241_, new_n_n234_, new_nxz160_f_,
    new_n_n222_, new_n_n219_, new_nmis11556_, new_n_n213_, new_n_n209_,
    new_nmis16748_, new_nmis16548_, new_nmis11593_, new_n_n185_,
    new_nmis16728_, new_n_n173_, new_n_n168_, new_nmis16596_, new_n_n154_,
    new_n_n146_, new_n_n139_, new_n_n129_, new_nmis16572_, new_nmis7564_,
    new_nmis15328_, new_nmis9061_, new_nmis15065_, new_n_n106_, new_n_n98_,
    new_n_n3_, new_n_n381_, new_n_n375_, new_n_n351_, new_n_n345_,
    new_n_n339_, new_n_n333_, new_n_n327_, new_n_n321_, new_ncomppar_p_,
    new_nrxz0_p_, new_naxz1_p_, new_n_n293_, new_n_n287_, new_n_n281_,
    new_n_n275_, new_n_n269_, new_n_n264_, new_n_n257_, new_ntxwrd7_p_,
    new_n_n240_, new_n_n235_, new_n_n229_, new_n_n223_, new_n_n218_,
    new_nmis11565_, new_nmis10130_, new_nmis8641_, new_n_n204_,
    new_nmis15843_, new_nmis11594_, new_n_n186_, new_n_n181_, new_n_n174_,
    new_n_n167_, new_n_n160_, new_nmis16734_, new_n_n147_, new_nmis11550_,
    new_nmis16883_, new_n_n125_, new_nmis16752_, new_nmis16765_,
    new_n_n112_, new_nmis15062_, new_nmis16611_, new_n_n99_, new_n_n4_,
    new_nmis16746_, new_nmis16873_, new_n_n72_, new_n_n61_, new_n_n50_,
    new_nmis12425_, new_n_n76_, new_nmis16767_, new_n_n60_, new_n_n51_,
    new_nmis16657_, new_n_n75_, new_n_n70_, new_n_n63_, new_n_n52_,
    new_nmis16675_, new_nmis15855_, new_n_n71_, new_n_n62_, new_n_n53_,
    new_n_n0_, new_nmis16673_, new_n_n43_, new_n_n32_, new_n_n21_,
    new_n_n10_, new_nmis16646_, new_n_n42_, new_n_n33_, new_n_n20_,
    new_n_n11_, new_n_n41_, new_n_n30_, new_n_n23_, new_n_n12_, new_n_n40_,
    new_n_n31_, new_n_n22_, new_n_n13_, new_n_n69_, new_n_n58_, new_n_n47_,
    new_n_n36_, new_n_n25_, new_n_n14_, new_n_n68_, new_n_n59_, new_n_n46_,
    new_n_n37_, new_n_n24_, new_n_n15_, new_nmis16719_, new_nmis16023_,
    new_n_n45_, new_n_n34_, new_n_n27_, new_n_n16_, new_n_n80_,
    new_nmis15854_, new_n_n44_, new_n_n35_, new_n_n26_, new_n_n17_,
    new_nmis16792_, new_n_n79_, new_nmis16027_, new_n_n65_, new_n_n54_,
    new_n_n29_, new_n_n18_, new_nmis16895_, new_nmis16871_, new_n_n74_,
    new_n_n64_, new_n_n55_, new_n_n28_, new_n_n19_, new_n_n81_, new_n_n78_,
    new_nmis16750_, new_n_n67_, new_n_n56_, new_n_n49_, new_n_n38_,
    new_n_n82_, new_n_n77_, new_n_n73_, new_n_n66_, new_n_n57_, new_n_n48_,
    new_n_n39_;
  assign new_ntxwrd3_ = txwrd3;
  assign new_na_ = a;
  assign i1zzz0_p = new_ni1zzz0_p_;
  assign new_nqpr4_ = qpr4;
  assign new_ntxwrd2_ = txwrd2;
  assign new_nb_ = b;
  assign new_ni1zzz0_ = i1zzz0;
  assign new_ntxwrd5_ = txwrd5;
  assign v1zzz0_p = new_nv1zzz0_p_;
  assign new_nc_ = c;
  assign new_np1zzz0_ = p1zzz0;
  assign new_ntxwrd4_ = txwrd4;
  assign new_nxzfs_ = xzfs;
  assign new_ni1zzz2_ = i1zzz2;
  assign i1zzz3_p = new_ni1zzz3_p_;
  assign new_ni2zzz1_ = i2zzz1;
  assign i2zzz2_p = new_ni2zzz2_p_;
  assign new_np1zzz1_ = p1zzz1;
  assign new_np2zzz0_ = p2zzz0;
  assign new_nqpr1_ = qpr1;
  assign txwrd8_p = new_ntxwrd8_p_;
  assign v1zzz2_p = new_nv1zzz2_p_;
  assign v2zzz1_p = new_nv2zzz1_p_;
  assign new_ni1zzz1_ = i1zzz1;
  assign i1zzz4_p = new_ni1zzz4_p_;
  assign new_ni2zzz0_ = i2zzz0;
  assign i2zzz3_p = new_ni2zzz3_p_;
  assign new_np1zzz2_ = p1zzz2;
  assign new_np2zzz1_ = p2zzz1;
  assign new_nqpr0_ = qpr0;
  assign stw_f = new_nstw_f_;
  assign txwrd9_p = new_ntxwrd9_p_;
  assign v1zzz1_p = new_nv1zzz1_p_;
  assign v2zzz0_p = new_nv2zzz0_p_;
  assign xz163_p = new_nxz163_p_;
  assign c_p = new_nc_p_;
  assign enwin_p = new_nenwin_p_;
  assign i1zzz1_p = new_ni1zzz1_p_;
  assign new_ni1zzz4_ = i1zzz4;
  assign i2zzz0_p = new_ni2zzz0_p_;
  assign new_ni2zzz3_ = i2zzz3;
  assign new_ninfin_ = infin;
  assign new_np1zzz3_ = p1zzz3;
  assign new_np2zzz2_ = p2zzz2;
  assign new_nqpr3_ = qpr3;
  assign new_ntxwrd1_ = txwrd1;
  assign txwrd6_p = new_ntxwrd6_p_;
  assign v1zzz4_p = new_nv1zzz4_p_;
  assign v2zzz3_p = new_nv2zzz3_p_;
  assign new_nvybb1_ = vybb1;
  assign i1zzz2_p = new_ni1zzz2_p_;
  assign new_ni1zzz3_ = i1zzz3;
  assign i2zzz1_p = new_ni2zzz1_p_;
  assign new_ni2zzz2_ = i2zzz2;
  assign new_np1zzz4_ = p1zzz4;
  assign new_np2zzz3_ = p2zzz3;
  assign new_nqpr2_ = qpr2;
  assign new_ntxwrd0_ = txwrd0;
  assign txwrd7_p = new_ntxwrd7_p_;
  assign v1zzz3_p = new_nv1zzz3_p_;
  assign v2zzz2_p = new_nv2zzz2_p_;
  assign new_nvybb0_ = vybb0;
  assign new_ncomppar_ = comppar;
  assign p1zzz4_p = new_np1zzz4_p_;
  assign p2zzz3_p = new_np2zzz3_p_;
  assign new_npsrw_ = psrw;
  assign xz162_p = new_nxz162_p_;
  assign new_nxz323_ = xz323;
  assign b_p = new_nb_p_;
  assign new_ncbt2_ = cbt2;
  assign new_nmmerr_ = mmerr;
  assign p1zzz3_p = new_np1zzz3_p_;
  assign p2zzz2_p = new_np2zzz2_p_;
  assign new_nryz_ = ryz;
  assign new_nxz324_ = xz324;
  assign p1zzz2_p = new_np1zzz2_p_;
  assign p2zzz1_p = new_np2zzz1_p_;
  assign xzfr1_p = new_nxzfr1_p_;
  assign new_nesrsum_ = esrsum;
  assign p1zzz1_p = new_np1zzz1_p_;
  assign p2zzz0_p = new_np2zzz0_p_;
  assign txwrd14_p = new_ntxwrd14_p_;
  assign xz161_p = new_nxz161_p_;
  assign a_p = new_na_p_;
  assign p1zzz0_p = new_np1zzz0_p_;
  assign new_nv1zzz7_ = v1zzz7;
  assign new_nv2zzz6_ = v2zzz6;
  assign new_nxz161_ = xz161;
  assign new_npfin_ = pfin;
  assign new_nstw_n_ = stw_n;
  assign new_nv2zzz7_ = v2zzz7;
  assign new_nvzzze_ = vzzze;
  assign new_nxz162_ = xz162;
  assign new_nxz320_ = xz320;
  assign axz0_p = new_naxz0_p_;
  assign new_ncbt1_ = cbt1;
  assign new_nslad0_ = slad0;
  assign txwrd15_p = new_ntxwrd15_p_;
  assign new_nv1zzz5_ = v1zzz5;
  assign new_nv2zzz4_ = v2zzz4;
  assign new_nxz163_ = xz163;
  assign new_nxz321_ = xz321;
  assign axz1_p = new_naxz1_p_;
  assign new_ncbt0_ = cbt0;
  assign new_nslad1_ = slad1;
  assign td_p = new_ntd_p_;
  assign new_nv1zzz6_ = v1zzz6;
  assign new_nv2zzz5_ = v2zzz5;
  assign new_nxz322_ = xz322;
  assign fsesr_p = new_nfsesr_p_;
  assign new_npybb5_ = pybb5;
  assign new_nslad2_ = slad2;
  assign new_ntxwrd14_ = txwrd14;
  assign new_nv1zzz3_ = v1zzz3;
  assign new_nv2zzz2_ = v2zzz2;
  assign new_nxz160_n_ = xz160_n;
  assign new_npybb4_ = pybb4;
  assign rptwin_p = new_nrptwin_p_;
  assign new_nslad3_ = slad3;
  assign txwrd12_p = new_ntxwrd12_p_;
  assign new_ntxwrd13_ = txwrd13;
  assign new_nv1zzz4_ = v1zzz4;
  assign new_nv2zzz3_ = v2zzz3;
  assign new_niclr_ = iclr;
  assign new_npybb3_ = pybb3;
  assign new_nrptwin_ = rptwin;
  assign txwrd11_p = new_ntxwrd11_p_;
  assign new_ntxwrd12_ = txwrd12;
  assign new_nv1zzz1_ = v1zzz1;
  assign new_nv2zzz0_ = v2zzz0;
  assign xz322_p = new_nxz322_p_;
  assign new_npybb2_ = pybb2;
  assign new_ntxwrd11_ = txwrd11;
  assign new_nv1zzz2_ = v1zzz2;
  assign new_nv2zzz1_ = v2zzz1;
  assign new_naxz1_ = axz1;
  assign new_ninzzze_ = inzzze;
  assign p2zzz7_p = new_np2zzz7_p_;
  assign txwrd13_p = new_ntxwrd13_p_;
  assign xz324_p = new_nxz324_p_;
  assign xzfs_p = new_nxzfs_p_;
  assign new_naxz0_ = axz0;
  assign p1zzz7_p = new_np1zzz7_p_;
  assign p2zzz6_p = new_np2zzz6_p_;
  assign new_npybb8_ = pybb8;
  assign new_nv1zzz0_ = v1zzz0;
  assign xzfr0_p = new_nxzfr0_p_;
  assign new_ninybb8_ = inybb8;
  assign p1zzz6_p = new_np1zzz6_p_;
  assign p2zzz5_p = new_np2zzz5_p_;
  assign new_npybb7_ = pybb7;
  assign rxz1_p = new_nrxz1_p_;
  assign new_nxzfr0_ = xzfr0;
  assign comppar_p = new_ncomppar_p_;
  assign new_nenwin_ = enwin;
  assign new_nofs1_ = ofs1;
  assign ofs2_p = new_nofs2_p_;
  assign p1zzz5_p = new_np1zzz5_p_;
  assign p2zzz4_p = new_np2zzz4_p_;
  assign new_npybb6_ = pybb6;
  assign new_npzzze_ = pzzze;
  assign rxz0_p = new_nrxz0_p_;
  assign new_ntxmess_n_ = txmess_n;
  assign new_ntxwrd15_ = txwrd15;
  assign xz323_p = new_nxz323_p_;
  assign new_nxzfr1_ = xzfr1;
  assign new_ni1zzz6_ = i1zzz6;
  assign i1zzz7_p = new_ni1zzz7_p_;
  assign new_ni2zzz5_ = i2zzz5;
  assign i2zzz6_p = new_ni2zzz6_p_;
  assign new_ninybb6_ = inybb6;
  assign ofs1_p = new_nofs1_p_;
  assign new_nofs2_ = ofs2;
  assign new_np1zzz5_ = p1zzz5;
  assign new_np2zzz4_ = p2zzz4;
  assign new_nrxz0_ = rxz0;
  assign ryz_p = new_nryz_p_;
  assign sbuff = new_nsbuff_;
  assign txwrd4_p = new_ntxwrd4_p_;
  assign v1zzz6_p = new_nv1zzz6_p_;
  assign v2zzz5_p = new_nv2zzz5_p_;
  assign xz160_f = new_nxz160_f_;
  assign xz320_p = new_nxz320_p_;
  assign new_ni1zzz5_ = i1zzz5;
  assign new_ni2zzz4_ = i2zzz4;
  assign i2zzz7_p = new_ni2zzz7_p_;
  assign new_ninybb7_ = inybb7;
  assign new_np1zzz6_ = p1zzz6;
  assign new_np2zzz5_ = p2zzz5;
  assign new_nrpten_ = rpten;
  assign new_nrxz1_ = rxz1;
  assign txwrd5_p = new_ntxwrd5_p_;
  assign v1zzz5_p = new_nv1zzz5_p_;
  assign v2zzz4_p = new_nv2zzz4_p_;
  assign i1zzz5_p = new_ni1zzz5_p_;
  assign i2zzz4_p = new_ni2zzz4_p_;
  assign new_ni2zzz7_ = i2zzz7;
  assign new_ninybb4_ = inybb4;
  assign new_np1zzz7_ = p1zzz7;
  assign new_np2zzz6_ = p2zzz6;
  assign qpr4_p = new_nqpr4_p_;
  assign txwrd2_p = new_ntxwrd2_p_;
  assign v2zzz7_p = new_nv2zzz7_p_;
  assign i1zzz6_p = new_ni1zzz6_p_;
  assign new_ni1zzz7_ = i1zzz7;
  assign i2zzz5_p = new_ni2zzz5_p_;
  assign new_ni2zzz6_ = i2zzz6;
  assign new_ninybb5_ = inybb5;
  assign new_np2zzz7_ = p2zzz7;
  assign txwrd3_p = new_ntxwrd3_p_;
  assign v1zzz7_p = new_nv1zzz7_p_;
  assign v2zzz6_p = new_nv2zzz6_p_;
  assign new_ninybb2_ = inybb2;
  assign new_npybb1_ = pybb1;
  assign qpr2_p = new_nqpr2_p_;
  assign txwrd0_p = new_ntxwrd0_p_;
  assign new_ntxwrd7_ = txwrd7;
  assign new_ntxwrd10_ = txwrd10;
  assign new_ninybb3_ = inybb3;
  assign new_npybb0_ = pybb0;
  assign qpr3_p = new_nqpr3_p_;
  assign txwrd1_p = new_ntxwrd1_p_;
  assign new_ntxwrd6_ = txwrd6;
  assign xz321_p = new_nxz321_p_;
  assign new_ninybb0_ = inybb0;
  assign qpr0_p = new_nqpr0_p_;
  assign new_ntxwrd9_ = txwrd9;
  assign new_ninybb1_ = inybb1;
  assign new_npsync_ = psync;
  assign qpr1_p = new_nqpr1_p_;
  assign txmess_f = new_ntxmess_f_;
  assign new_ntxwrd8_ = txwrd8;
  assign txwrd10_p = new_ntxwrd10_p_;
  assign new_nvfin_ = vfin;
  assign new_nsbuff_ = new_nrptwin_ | new_n_n30_;
  assign new_n_n378_ = new_nmis11587_ & new_np1zzz1_;
  assign new_np1zzz5_p_ = new_n_n369_ | new_n_n370_;
  assign new_n_n363_ = new_nmis11586_ & new_npybb1_;
  assign new_n_n356_ = new_nmis11585_ & new_np2zzz4_;
  assign new_ni1zzz0_p_ = new_n_n347_ | new_n_n348_;
  assign new_n_n341_ = new_nmis11582_ & new_ninybb4_;
  assign new_n_n334_ = new_nmis11581_ & new_ni1zzz7_;
  assign new_ni2zzz3_p_ = new_n_n325_ | new_n_n326_;
  assign new_n_n319_ = new_nmis11584_ & new_ninybb7_;
  assign new_nxzfr1_p_ = new_n_n313_ | new_n_n314_;
  assign new_nofs1_p_ = new_n_n22_ & new_npsync_;
  assign new_n_n304_ = new_nmis15843_ & new_n_n41_;
  assign new_n_n298_ = new_nmis11589_ & new_nv1zzz0_;
  assign new_nv1zzz4_p_ = new_n_n289_ | new_n_n290_;
  assign new_n_n283_ = new_nmis11590_ & new_nvybb1_;
  assign new_n_n276_ = new_nmis11591_ & new_nv2zzz3_;
  assign new_nv2zzz7_p_ = new_n_n267_ | new_n_n268_;
  assign new_n_n262_ = new_ni1zzz3_ & new_nmis11594_;
  assign new_ntxwrd6_p_ = new_n_n253_ | new_n_n252_ | new_n_n251_;
  assign new_n_n246_ = new_nmis16627_ & new_nmis11593_;
  assign new_nxz323_p_ = new_n_n232_ | new_n_n233_;
  assign new_n_n226_ = new_n_n56_ & new_n_n21_ & new_nmis15083_;
  assign new_nmis16706_ = new_n_n220_ | new_n_n219_ | new_n_n218_;
  assign new_nmis11584_ = new_n_n5_ & new_n_n19_;
  assign new_n_n212_ = new_nmis11560_ & new_nmis8027_;
  assign new_nmis16544_ = new_n_n207_ | new_nxz320_p_;
  assign new_n_n201_ = new_nmis9174_ & new_nc_;
  assign new_n_n197_ = new_nmis16555_ & new_naxz1_;
  assign new_n_n178_ = new_nv1zzz5_ & new_nvfin_;
  assign new_nmis16631_ = new_n_n169_ | new_n_n168_ | new_n_n167_;
  assign new_n_n161_ = new_nmis11547_ & new_nmis16611_;
  assign new_n_n153_ = new_nv2zzz5_ & new_nvfin_;
  assign new_nmis11560_ = new_n_n22_ & new_n_n36_;
  assign new_nmis10125_ = new_nmis7564_ | new_nxz160_n_;
  assign new_nmis16690_ = new_n_n134_ | new_n_n135_;
  assign new_nmis9174_ = new_n_n113_ | new_nqpr3_ | new_ntxmess_n_ | new_nmis8768_;
  assign new_n_n109_ = new_nmis11549_ & new_ntxwrd1_;
  assign new_n_n105_ = new_nv2zzz2_ & new_nvfin_;
  assign new_nmis16742_ = new_n_n51_ | new_n_n50_;
  assign new_nmis9255_ = new_nc_ | new_nb_;
  assign new_nmis16866_ = new_n_n83_ | new_n_n84_;
  assign new_n_n371_ = new_nmis11588_ & new_npybb5_;
  assign new_n_n370_ = new_nmis11587_ & new_np1zzz5_;
  assign new_n_n364_ = new_nmis11585_ & new_np2zzz0_;
  assign new_n_n355_ = new_nmis11586_ & new_npybb5_;
  assign new_n_n349_ = new_nmis11586_ & new_npybb8_;
  assign new_ni1zzz4_p_ = new_n_n339_ | new_n_n340_;
  assign new_ni1zzz7_p_ = new_n_n333_ | new_n_n334_;
  assign new_n_n326_ = new_nmis11583_ & new_ni2zzz3_;
  assign new_n_n320_ = new_nmis11583_ & new_ni2zzz6_;
  assign new_n_n314_ = new_nmis16613_ & new_nxzfr1_;
  assign new_nofs2_p_ = new_nofs1_ & new_n_n22_;
  assign new_na_p_ = new_n_n19_ & new_nmis16748_;
  assign new_n_n297_ = new_nmis11590_ & new_nv1zzz1_;
  assign new_n_n291_ = new_nmis11590_ & new_nv1zzz4_;
  assign new_nv2zzz0_p_ = new_n_n281_ | new_n_n282_;
  assign new_nv2zzz3_p_ = new_n_n275_ | new_n_n276_;
  assign new_n_n268_ = new_nmis11591_ & new_nv2zzz7_;
  assign new_ntxwrd3_p_ = new_n_n262_ | new_n_n261_ | new_n_n260_;
  assign new_n_n253_ = new_ni1zzz6_ & new_nmis11594_;
  assign new_n_n247_ = new_ni2zzz1_ & new_nmis11594_;
  assign new_n_n233_ = new_nmis16730_ & new_nxz323_;
  assign new_n_n227_ = new_nmis9071_ & new_nxz161_;
  assign new_n_n220_ = new_n_n25_ & new_nmis16701_ & new_n_n30_;
  assign new_nmis11583_ = new_n_n19_ & new_nmis16887_;
  assign new_nmis8027_ = new_nxz161_ | new_nxz163_ | new_nmis7564_ | new_nxz162_ | new_n_n67_;
  assign new_n_n208_ = new_n_n66_ & new_nofs1_p_ & new_n_n68_ & new_nxzfs_ & new_n_n70_ & new_n_n65_;
  assign new_n_n200_ = new_n_n13_ & new_n_n14_;
  assign new_nmis16553_ = new_n_n196_ | new_n_n197_;
  assign new_nmis16726_ = new_n_n184_ | new_n_n183_ | new_n_n182_;
  assign new_n_n169_ = new_nv2zzz0_ & new_nvfin_;
  assign new_n_n162_ = new_nmis11546_ & new_np2zzz2_;
  assign new_n_n152_ = new_nmis11548_ & new_ntxwrd13_;
  assign new_n_n145_ = new_nmis11562_ & new_nv2zzz7_;
  assign new_nmis9071_ = new_n_n140_ | new_nxz320_p_;
  assign new_n_n136_ = new_nofs1_p_ & new_nxzfs_;
  assign new_n_n113_ = new_nmis16895_ & new_n_n42_;
  assign new_n_n110_ = new_nmis11548_ & new_ntxwrd0_;
  assign new_n_n104_ = new_nmis11548_ & new_ntxwrd10_;
  assign new_n_n97_ = new_nmis11549_ & new_ntxwrd13_;
  assign new_nmis16577_ = new_n_n89_ | new_n_n90_;
  assign new_n_n85_ = new_n_n70_ & new_n_n56_;
  assign new_n_n379_ = new_nmis11588_ & new_npybb1_;
  assign new_n_n372_ = new_nmis11587_ & new_np1zzz4_;
  assign new_np2zzz5_p_ = new_n_n353_ | new_n_n354_;
  assign new_n_n347_ = new_nmis11582_ & new_ninybb1_;
  assign new_ni1zzz3_p_ = new_n_n341_ | new_n_n342_;
  assign new_n_n335_ = new_nmis11582_ & new_ninybb7_;
  assign new_n_n325_ = new_nmis11584_ & new_ninybb4_;
  assign new_n_n318_ = new_nmis11583_ & new_ni2zzz7_;
  assign new_n_n316_ = new_nmis10130_ & new_nxzfr0_;
  assign new_n_n309_ = new_nrxz0_ & new_n_n33_ & new_nmis8641_;
  assign new_nv1zzz1_p_ = new_n_n295_ | new_n_n296_;
  assign new_n_n289_ = new_nmis11590_ & new_nv1zzz5_;
  assign new_nv1zzz7_p_ = new_n_n283_ | new_n_n284_;
  assign new_n_n277_ = new_nmis11592_ & new_nv2zzz3_;
  assign new_n_n267_ = new_nmis11592_ & new_nvybb1_;
  assign new_n_n260_ = new_nmis15080_ & new_nmis16726_;
  assign new_n_n255_ = new_np1zzz5_ & new_nmis15081_;
  assign new_ntxwrd9_p_ = new_n_n246_ | new_n_n247_;
  assign new_n_n232_ = new_n_n51_ & new_nmis15083_ & new_nmis11578_;
  assign new_n_n225_ = new_nxz162_ & new_nmis16588_;
  assign new_nmis16790_ = new_n_n221_ | new_nstw_n_;
  assign new_nmis11582_ = new_n_n4_ & new_n_n19_;
  assign new_nmis15083_ = new_nmis11560_ & new_nxz320_;
  assign new_nmis16541_ = new_n_n205_ | new_n_n206_;
  assign new_n_n202_ = new_n_n30_ & new_n_n12_ & new_n_n72_ & new_n_n11_ & new_n_n58_ & new_n_n42_;
  assign new_n_n198_ = new_n_n16_ & new_n_n61_;
  assign new_n_n184_ = new_nv1zzz3_ & new_nvfin_;
  assign new_n_n176_ = new_nmis11549_ & new_ntxwrd6_;
  assign new_nmis16609_ = new_n_n162_ | new_n_n161_ | new_n_n160_;
  assign new_n_n151_ = new_nmis11549_ & new_ntxwrd14_;
  assign new_n_n144_ = new_nmis11560_ & new_n_n20_;
  assign new_nmis16754_ = new_n_n141_ | new_nxz320_p_;
  assign new_n_n137_ = new_nenwin_ & new_n_n22_;
  assign new_n_n123_ = new_n_n53_ & new_n_n61_;
  assign new_n_n118_ = new_nmis16675_ & new_nmis15650_;
  assign new_n_n103_ = new_nmis11549_ & new_ntxwrd11_;
  assign new_nmis16778_ = new_n_n95_ | new_n_n96_;
  assign new_n_n92_ = new_naxz1_ & new_nmis16719_;
  assign new_n_n86_ = new_nslad1_ & new_nxz161_;
  assign new_nstw_f_ = new_n_n383_ | new_nryz_;
  assign new_np1zzz1_p_ = new_n_n377_ | new_n_n378_;
  assign new_np1zzz4_p_ = new_n_n371_ | new_n_n372_;
  assign new_n_n354_ = new_nmis11585_ & new_np2zzz5_;
  assign new_n_n348_ = new_nmis11581_ & new_ni1zzz0_;
  assign new_n_n342_ = new_nmis11581_ & new_ni1zzz3_;
  assign new_n_n336_ = new_nmis11581_ & new_ni1zzz6_;
  assign new_ni2zzz4_p_ = new_n_n323_ | new_n_n324_;
  assign new_ni2zzz7_p_ = new_n_n317_ | new_n_n318_;
  assign new_n_n315_ = new_n_n7_ & new_n_n0_ & new_nmis15083_;
  assign new_n_n310_ = new_nmis16541_ & new_nrxz1_;
  assign new_n_n296_ = new_nmis11589_ & new_nv1zzz1_;
  assign new_n_n290_ = new_nmis11589_ & new_nv1zzz4_;
  assign new_n_n284_ = new_nmis11589_ & new_nv1zzz7_;
  assign new_n_n278_ = new_nmis11591_ & new_nv2zzz2_;
  assign new_ntxwrd0_p_ = new_n_n19_ & new_nmis16591_;
  assign new_n_n261_ = new_np1zzz3_ & new_nmis15081_;
  assign new_n_n254_ = new_nmis15080_ & new_nmis16732_;
  assign new_n_n248_ = new_nmis15080_ & new_nmis16631_;
  assign new_nxz324_p_ = new_n_n230_ | new_n_n231_;
  assign new_nxz162_p_ = new_n_n224_ | new_n_n225_;
  assign new_n_n221_ = new_nmis11556_ & new_na_;
  assign new_nmis11581_ = new_n_n19_ & new_nmis16891_;
  assign new_nmis16613_ = new_n_n211_ | new_nmis10130_;
  assign new_n_n207_ = new_nmis15964_ & new_n_n22_;
  assign new_nmis16762_ = new_n_n200_ | new_n_n201_;
  assign new_n_n199_ = new_nmis9061_ & new_naxz0_;
  assign new_n_n183_ = new_nmis11548_ & new_ntxwrd3_;
  assign new_n_n177_ = new_nmis11548_ & new_ntxwrd5_;
  assign new_n_n170_ = new_np1zzz7_ & new_nmis11546_;
  assign new_nmis16736_ = new_n_n150_ | new_n_n149_ | new_n_n148_;
  assign new_nmis15339_ = new_n_n144_ | new_nxz320_p_;
  assign new_n_n141_ = new_nmis11560_ & new_nmis7564_;
  assign new_nmis16786_ = new_n_n136_ | new_n_n137_;
  assign new_nmis16724_ = new_n_n33_ | new_n_n32_;
  assign new_n_n119_ = new_n_n36_ & new_nmis16673_;
  assign new_nmis16598_ = new_n_n102_ | new_n_n101_ | new_n_n100_;
  assign new_nmis16604_ = new_n_n56_ | new_n_n64_;
  assign new_n_n91_ = new_n_n54_ & new_naxz0_ & new_n_n53_;
  assign new_nmis16864_ = new_n_n85_ | new_n_n86_;
  assign new_n_n368_ = new_nmis11587_ & new_np1zzz6_;
  assign new_np2zzz2_p_ = new_n_n359_ | new_n_n360_;
  assign new_n_n344_ = new_nmis11581_ & new_ni1zzz2_;
  assign new_ni1zzz6_p_ = new_n_n335_ | new_n_n336_;
  assign new_nqpr0_p_ = new_n_n307_ | new_n_n308_;
  assign new_n_n301_ = new_nqpr3_ & new_nmis16548_ & new_n_n19_;
  assign new_nv2zzz2_p_ = new_n_n277_ | new_n_n278_;
  assign new_ntxwrd1_p_ = new_n_n265_ | new_n_n266_;
  assign new_ntxwrd13_p_ = new_n_n245_ | new_n_n244_ | new_n_n243_;
  assign new_nxz320_p_ = new_nmis11560_ & new_n_n57_;
  assign new_n_n211_ = new_nmis11560_ & new_n_n7_;
  assign new_n_n205_ = new_n_n22_ & new_n_n32_;
  assign new_nmis11591_ = new_n_n19_ & new_nmis16893_;
  assign new_n_n190_ = new_nmis15065_ & new_ntxwrd2_;
  assign new_n_n150_ = new_nv2zzz6_ & new_nvfin_;
  assign new_nmis16730_ = new_n_n143_ | new_nmis15339_;
  assign new_nmis16588_ = new_n_n139_ | new_nmis9071_;
  assign new_n_n133_ = new_na_ & new_nmis16716_;
  assign new_nmis11154_ = new_n_n127_ | new_n_n128_;
  assign new_n_n102_ = new_nv2zzz3_ & new_nvfin_;
  assign new_n_n95_ = new_nslad3_ & new_n_n52_;
  assign new_nmis16579_ = new_n_n87_ | new_n_n88_;
  assign new_nmis16670_ = new_n_n64_ | new_nmis15854_ | new_n_n57_;
  assign new_n_n9_ = ~new_nofs1_;
  assign new_n_n367_ = new_nmis11588_ & new_npybb7_;
  assign new_n_n361_ = new_nmis11586_ & new_npybb2_;
  assign new_n_n343_ = new_nmis11582_ & new_ninybb3_;
  assign new_n_n337_ = new_nmis11582_ & new_ninybb6_;
  assign new_n_n308_ = new_n_n15_ & new_n_n52_;
  assign new_n_n302_ = new_nqpr2_ & new_n_n58_ & new_nmis15843_;
  assign new_n_n285_ = new_nmis11590_ & new_nv1zzz7_;
  assign new_ntxwrd4_p_ = new_n_n259_ | new_n_n258_ | new_n_n257_;
  assign new_n_n245_ = new_np2zzz5_ & new_nmis15081_;
  assign new_n_n238_ = new_nmis16583_ & new_nmis11593_;
  assign new_nmis16879_ = new_n_n210_ | new_nofs1_p_;
  assign new_n_n206_ = new_nmis16544_ & new_n_n25_;
  assign new_nmis11592_ = new_n_n18_ & new_n_n19_;
  assign new_n_n191_ = new_nmis15062_ & new_ntxwrd1_;
  assign new_n_n149_ = new_nmis11548_ & new_ntxwrd14_;
  assign new_nmis11578_ = new_nxz322_ & new_nxz321_;
  assign new_nmis16701_ = new_n_n132_ | new_n_n133_;
  assign new_n_n132_ = new_nmis9255_ & new_ntxwrd0_ & new_nmis7401_;
  assign new_nmis16887_ = new_n_n29_ | new_n_n28_;
  assign new_n_n101_ = new_nmis11548_ & new_ntxwrd11_;
  assign new_n_n96_ = new_nslad2_ & new_nqpr0_;
  assign new_n_n88_ = new_naxz0_ & new_nmmerr_;
  assign new_nmis16665_ = new_n_n63_ | new_nmis15855_ | new_n_n57_;
  assign new_n_n369_ = new_nmis11588_ & new_npybb6_;
  assign new_n_n362_ = new_nmis11585_ & new_np2zzz1_;
  assign new_n_n357_ = new_nmis11586_ & new_npybb4_;
  assign new_n_n350_ = new_nmis11585_ & new_np2zzz7_;
  assign new_nb_p_ = new_n_n19_ & new_nmis16760_;
  assign new_nqpr3_p_ = new_n_n301_ | new_n_n302_;
  assign new_n_n292_ = new_nmis11589_ & new_nv1zzz3_;
  assign new_n_n252_ = new_np1zzz6_ & new_nmis15081_;
  assign new_ntxwrd11_p_ = new_n_n19_ & new_nmis16596_;
  assign new_n_n239_ = new_ni2zzz7_ & new_nmis11594_;
  assign new_nmis16629_ = new_nmis11565_ | new_n_n52_;
  assign new_nmis11589_ = new_n_n19_ & new_nmis16889_;
  assign new_n_n192_ = new_np1zzz1_ & new_npfin_;
  assign new_n_n148_ = new_nmis11549_ & new_ntxwrd15_;
  assign new_n_n140_ = new_nmis11560_ & new_nmis10125_;
  assign new_n_n134_ = new_n_n23_ & new_nqpr2_ & new_nmis16780_;
  assign new_n_n100_ = new_nmis11549_ & new_ntxwrd12_;
  assign new_n_n94_ = new_nqpr0_ & new_nslad0_;
  assign new_n_n90_ = new_naxz0_ & new_n_n54_;
  assign new_n_n83_ = new_n_n68_ & new_nxz160_n_;
  assign new_np1zzz6_p_ = new_n_n367_ | new_n_n368_;
  assign new_np2zzz1_p_ = new_n_n361_ | new_n_n362_;
  assign new_np2zzz4_p_ = new_n_n355_ | new_n_n356_;
  assign new_np2zzz7_p_ = new_n_n349_ | new_n_n350_;
  assign new_nc_p_ = new_n_n19_ & new_nmis16762_;
  assign new_n_n303_ = new_nqpr2_ & new_nmis16581_ & new_n_n19_;
  assign new_nv1zzz0_p_ = new_n_n297_ | new_n_n298_;
  assign new_ntxwrd10_p_ = new_nmis16609_ & new_n_n19_;
  assign new_ntxwrd12_p_ = new_n_n19_ & new_nmis16623_;
  assign new_ntxwrd15_p_ = new_n_n238_ | new_n_n239_;
  assign new_nmis16581_ = new_nmis16629_ | new_n_n23_;
  assign new_n_n196_ = new_n_n16_ & new_naxz0_ & new_n_n53_;
  assign new_nmis11590_ = new_n_n17_ & new_n_n19_;
  assign new_n_n143_ = new_nmis11560_ & new_n_n50_;
  assign new_nmis15848_ = new_nxz320_ & new_nxz161_ & new_n_n21_;
  assign new_n_n135_ = new_nqpr1_ & new_n_n41_ & new_nmis16778_;
  assign new_nmis16625_ = new_n_n99_ | new_n_n98_ | new_n_n97_;
  assign new_nmis16780_ = new_n_n93_ | new_n_n94_;
  assign new_n_n89_ = new_naxz1_ & new_nesrsum_;
  assign new_n_n84_ = new_nslad0_ & new_n_n67_;
  assign new_ntd_p_ = new_n_n19_ & new_nmis16706_;
  assign new_n_n376_ = new_nmis11587_ & new_np1zzz2_;
  assign new_n_n365_ = new_nmis11588_ & new_npybb8_;
  assign new_n_n358_ = new_nmis11585_ & new_np2zzz3_;
  assign new_n_n317_ = new_nmis11584_ & new_ninybb8_;
  assign new_nxzfs_p_ = new_npsrw_ & new_nmis16879_ & new_nmis16788_;
  assign new_n_n306_ = new_nqpr0_ & new_n_n23_ & new_n_n15_;
  assign new_naxz0_p_ = new_n_n19_ & new_nmis16615_;
  assign new_nv1zzz3_p_ = new_n_n291_ | new_n_n292_;
  assign new_n_n251_ = new_nmis15080_ & new_nmis16633_;
  assign new_ntxwrd14_p_ = new_n_n242_ | new_n_n241_ | new_n_n240_;
  assign new_nxz322_p_ = new_n_n234_ | new_n_n235_;
  assign new_n_n228_ = new_n_n21_ & new_nmis15083_;
  assign new_nmis11547_ = new_n_n46_ & new_n_n47_;
  assign new_n_n194_ = new_nmis16593_ & new_nmis11547_;
  assign new_n_n187_ = new_nmis15062_ & new_ntxwrd2_;
  assign new_n_n180_ = new_nmis11548_ & new_ntxwrd4_;
  assign new_n_n172_ = new_nmis16620_ & new_nmis11547_;
  assign new_n_n163_ = new_nmis11562_ & new_nv2zzz1_;
  assign new_nmis16712_ = new_n_n129_ | new_n_n130_;
  assign new_n_n126_ = new_ncomppar_ & new_nmis16579_;
  assign new_nmis15964_ = new_n_n119_ | new_n_n118_ | new_n_n121_ | new_n_n120_ | new_n_n116_ | new_n_n122_ | new_n_n117_;
  assign new_nmis8768_ = new_n_n52_ | new_nqpr1_ | new_n_n41_;
  assign new_nmis16593_ = new_n_n111_ | new_n_n110_ | new_n_n109_;
  assign new_n_n107_ = new_nmis11548_ & new_ntxwrd7_;
  assign new_n_n5_ = ~new_nmis16887_;
  assign new_nfsesr_p_ = new_n_n381_ | new_n_n382_;
  assign new_np1zzz2_p_ = new_n_n375_ | new_n_n376_;
  assign new_np2zzz0_p_ = new_n_n363_ | new_n_n364_;
  assign new_np2zzz3_p_ = new_n_n357_ | new_n_n358_;
  assign new_ntxmess_f_ = new_nmis11565_ | new_nryz_;
  assign new_n_n313_ = new_nxzfr0_ & new_nmis15083_ & new_n_n0_ & new_n_n1_;
  assign new_n_n305_ = new_nqpr1_ & new_nmis16629_ & new_n_n19_;
  assign new_n_n299_ = new_nqpr2_ & new_n_n42_ & new_nmis15843_ & new_nqpr3_;
  assign new_n_n286_ = new_nmis11589_ & new_nv1zzz6_;
  assign new_n_n259_ = new_ni1zzz4_ & new_nmis11594_;
  assign new_n_n242_ = new_np2zzz6_ & new_nmis15081_;
  assign new_n_n236_ = new_nxz320_p_ & new_nxz321_;
  assign new_nxz161_p_ = new_n_n226_ | new_n_n227_;
  assign new_nenwin_p_ = new_npsrw_ & new_nmis16786_ & new_nmis16788_;
  assign new_n_n193_ = new_np1zzz0_ & new_nmis11546_;
  assign new_n_n188_ = new_np1zzz2_ & new_npfin_;
  assign new_n_n179_ = new_nmis11549_ & new_ntxwrd5_;
  assign new_nmis16618_ = new_n_n172_ | new_n_n171_ | new_n_n170_;
  assign new_n_n156_ = new_nmis11546_ & new_np2zzz4_;
  assign new_n_n130_ = new_nesrsum_ & new_n_n32_ & new_nrxz1_;
  assign new_nmis16565_ = new_nmis11556_ | new_n_n126_ | new_n_n125_;
  assign new_n_n122_ = new_nslad2_ & new_nmis16670_;
  assign new_n_n115_ = new_n_n39_ & new_n_n40_;
  assign new_n_n111_ = new_nv1zzz0_ & new_nvfin_;
  assign new_n_n108_ = new_nv1zzz7_ & new_nvfin_;
  assign new_n_n6_ = ~new_nmis15650_;
  assign new_n_n377_ = new_nmis11588_ & new_npybb2_;
  assign new_np1zzz7_p_ = new_n_n365_ | new_n_n366_;
  assign new_n_n359_ = new_nmis11586_ & new_npybb3_;
  assign new_ni2zzz1_p_ = new_n_n329_ | new_n_n330_;
  assign new_n_n323_ = new_nmis11584_ & new_ninybb5_;
  assign new_n_n307_ = new_n_n19_ & new_nqpr0_ & new_nmis11565_;
  assign new_n_n300_ = new_nmis16546_ & new_nqpr4_ & new_n_n19_;
  assign new_n_n279_ = new_nmis11592_ & new_nv2zzz2_;
  assign new_n_n266_ = new_ni1zzz1_ & new_nmis11594_;
  assign new_n_n244_ = new_ni2zzz5_ & new_nmis11594_;
  assign new_n_n237_ = new_nmis15083_ & new_n_n20_;
  assign new_nmis11585_ = new_n_n19_ & new_nmis16885_;
  assign new_n_n215_ = new_nmis11154_ & new_n_n30_ & new_n_n62_ & new_nmis7401_;
  assign new_nmis16591_ = new_n_n195_ | new_n_n194_ | new_n_n193_;
  assign new_nmis16585_ = new_n_n185_ | new_n_n187_ | new_n_n186_ | new_n_n188_;
  assign new_nmis16732_ = new_n_n178_ | new_n_n177_ | new_n_n176_;
  assign new_n_n165_ = new_nmis15062_ & new_ntxwrd9_;
  assign new_nmis16623_ = new_n_n156_ | new_n_n155_ | new_n_n154_;
  assign new_nmis16710_ = new_n_n131_ | new_n_n24_;
  assign new_n_n127_ = new_n_n60_ & new_n_n42_ & new_nmis16690_ & new_n_n58_;
  assign new_n_n121_ = new_nmis16646_ & new_nslad1_;
  assign new_n_n114_ = new_n_n58_ & new_nmis15328_;
  assign new_nmis16893_ = new_n_n45_ | new_n_n44_;
  assign new_nmis16620_ = new_n_n108_ | new_n_n107_ | new_n_n106_;
  assign new_n_n7_ = ~new_nxzfr0_;
  assign new_n_n383_ = new_n_n49_ & new_nmis11547_ & new_nmis16790_;
  assign new_n_n366_ = new_nmis11587_ & new_np1zzz7_;
  assign new_n_n360_ = new_nmis11585_ & new_np2zzz2_;
  assign new_n_n330_ = new_nmis11583_ & new_ni2zzz1_;
  assign new_n_n324_ = new_nmis11583_ & new_ni2zzz4_;
  assign new_nqpr1_p_ = new_n_n305_ | new_n_n306_;
  assign new_nqpr4_p_ = new_n_n299_ | new_n_n300_;
  assign new_nv2zzz5_p_ = new_n_n271_ | new_n_n272_;
  assign new_n_n272_ = new_nmis11591_ & new_nv2zzz5_;
  assign new_n_n243_ = new_nmis15080_ & new_nmis16734_;
  assign new_nxz321_p_ = new_n_n236_ | new_n_n237_;
  assign new_nmis11586_ = new_n_n3_ & new_n_n19_;
  assign new_n_n216_ = new_ncomppar_ & new_nmis16572_;
  assign new_n_n195_ = new_ni1zzz0_ & new_ninfin_;
  assign new_n_n189_ = new_nmis11562_ & new_nv1zzz1_;
  assign new_n_n171_ = new_ni1zzz7_ & new_ninfin_;
  assign new_n_n164_ = new_nmis15065_ & new_ntxwrd10_;
  assign new_n_n157_ = new_ni2zzz3_ & new_ninfin_;
  assign new_n_n131_ = new_n_n25_ & new_n_n60_ & new_nmis7401_;
  assign new_n_n128_ = new_ntxwrd0_ & new_nmis9255_;
  assign new_n_n120_ = new_nslad3_ & new_nmis16665_;
  assign new_nmis16758_ = new_n_n114_ | new_nmis8768_ | new_nqpr4_ | new_ntxmess_n_;
  assign new_nmis11546_ = new_n_n46_ & new_npfin_;
  assign new_nmis11549_ = new_n_n48_ & new_n_n49_;
  assign new_n_n8_ = ~new_nofs2_;
  assign new_np1zzz0_p_ = new_n_n379_ | new_n_n380_;
  assign new_n_n373_ = new_nmis11588_ & new_npybb4_;
  assign new_n_n353_ = new_nmis11586_ & new_npybb6_;
  assign new_n_n346_ = new_nmis11581_ & new_ni1zzz1_;
  assign new_ni1zzz5_p_ = new_n_n337_ | new_n_n338_;
  assign new_n_n331_ = new_nmis11584_ & new_ninybb1_;
  assign new_n_n329_ = new_nmis11584_ & new_ninybb2_;
  assign new_n_n322_ = new_nmis11583_ & new_ni2zzz5_;
  assign new_nrptwin_p_ = new_n_n19_ & new_nmis16722_;
  assign new_nrxz1_p_ = new_n_n309_ | new_n_n310_;
  assign new_n_n295_ = new_nmis11590_ & new_nv1zzz2_;
  assign new_n_n288_ = new_nmis11589_ & new_nv1zzz5_;
  assign new_nv2zzz1_p_ = new_n_n279_ | new_n_n280_;
  assign new_n_n273_ = new_nmis11592_ & new_nv2zzz5_;
  assign new_n_n271_ = new_nmis11592_ & new_nv2zzz6_;
  assign new_ntxwrd2_p_ = new_n_n263_ | new_n_n264_;
  assign new_ntxwrd5_p_ = new_n_n256_ | new_n_n255_ | new_n_n254_;
  assign new_n_n249_ = new_np2zzz0_ & new_nmis15081_;
  assign new_n_n231_ = new_nmis16740_ & new_nxz324_;
  assign new_nxz163_p_ = new_n_n222_ | new_n_n223_;
  assign new_nmis11587_ = new_n_n19_ & new_nmis16883_;
  assign new_n_n217_ = new_na_ & new_nmis16565_;
  assign new_nmis16722_ = new_nmis15847_ | new_n_n214_ | new_n_n213_;
  assign new_nmis16788_ = new_n_n9_ | new_n_n8_;
  assign new_nmis16760_ = new_n_n202_ | new_n_n203_;
  assign new_nmis16615_ = new_n_n198_ | new_n_n199_;
  assign new_nmis16606_ = new_n_n189_ | new_n_n191_ | new_n_n190_ | new_n_n192_;
  assign new_n_n182_ = new_nmis11549_ & new_ntxwrd4_;
  assign new_n_n175_ = new_nv1zzz6_ & new_nvfin_;
  assign new_nmis16627_ = new_n_n163_ | new_n_n165_ | new_n_n164_ | new_n_n166_;
  assign new_n_n158_ = new_nmis16598_ & new_nmis11547_;
  assign new_nmis16583_ = new_n_n147_ | new_n_n146_ | new_n_n145_;
  assign new_nmis16740_ = new_n_n142_ | new_nmis15339_;
  assign new_n_n138_ = new_nmis16604_ & new_nmis11560_;
  assign new_nmis16885_ = new_n_n27_ | new_n_n26_;
  assign new_nmis7401_ = new_n_n123_ | new_n_n43_;
  assign new_nmis15650_ = new_n_n37_ | new_nslad3_ | new_n_n36_ | new_nslad2_;
  assign new_n_n116_ = new_nmis12425_ & new_n_n37_;
  assign new_nmis16555_ = new_n_n61_ | new_nmis9061_;
  assign new_nmis11548_ = new_nmis16792_ & new_n_n49_;
  assign new_n_n93_ = new_n_n52_ & new_nslad1_;
  assign new_nmis16858_ = new_nmis16873_ & new_nmis16871_;
  assign new_n_n1_ = ~new_nxzfr1_;
  assign new_n_n380_ = new_nmis11587_ & new_np1zzz0_;
  assign new_n_n374_ = new_nmis11587_ & new_np1zzz3_;
  assign new_np2zzz6_p_ = new_n_n351_ | new_n_n352_;
  assign new_ni1zzz1_p_ = new_n_n345_ | new_n_n346_;
  assign new_n_n338_ = new_nmis11581_ & new_ni1zzz5_;
  assign new_n_n332_ = new_nmis11583_ & new_ni2zzz0_;
  assign new_ni2zzz2_p_ = new_n_n327_ | new_n_n328_;
  assign new_ni2zzz5_p_ = new_n_n321_ | new_n_n322_;
  assign new_nxzfr0_p_ = new_n_n315_ | new_n_n316_;
  assign new_n_n311_ = new_n_n25_ & new_nrxz0_ & new_nmis16544_;
  assign new_nv1zzz2_p_ = new_n_n293_ | new_n_n294_;
  assign new_nv1zzz5_p_ = new_n_n287_ | new_n_n288_;
  assign new_n_n280_ = new_nmis11591_ & new_nv2zzz1_;
  assign new_n_n274_ = new_nmis11591_ & new_nv2zzz4_;
  assign new_nv2zzz6_p_ = new_n_n269_ | new_n_n270_;
  assign new_n_n265_ = new_nmis16606_ & new_nmis11593_;
  assign new_n_n256_ = new_ni1zzz5_ & new_nmis11594_;
  assign new_n_n250_ = new_ni2zzz0_ & new_nmis11594_;
  assign new_n_n230_ = new_n_n34_ & new_nmis11550_ & new_nmis11560_;
  assign new_n_n224_ = new_nmis15848_ & new_n_n64_ & new_nmis11560_;
  assign new_nmis11588_ = new_n_n2_ & new_n_n19_;
  assign new_nmis16569_ = new_n_n217_ | new_n_n216_ | new_n_n215_;
  assign new_n_n214_ = new_nmis16724_ & new_nrptwin_;
  assign new_n_n210_ = new_nxzfs_ & new_n_n22_;
  assign new_n_n203_ = new_nmis16758_ & new_nb_;
  assign new_nmis16546_ = new_nmis16548_ | new_n_n58_;
  assign new_nmis15081_ = new_nmis11593_ & new_npfin_;
  assign new_nmis15080_ = new_nmis11593_ & new_n_n47_;
  assign new_nmis16633_ = new_n_n175_ | new_n_n174_ | new_n_n173_;
  assign new_n_n166_ = new_np2zzz1_ & new_npfin_;
  assign new_n_n159_ = new_nmis11546_ & new_np2zzz3_;
  assign new_n_n155_ = new_nmis16625_ & new_nmis11547_;
  assign new_n_n142_ = new_nmis11560_ & new_nmis16742_;
  assign new_nmis16602_ = new_n_n138_ | new_nmis9071_;
  assign new_nmis16891_ = new_ninzzze_ | new_n_n28_;
  assign new_n_n124_ = new_nmis7401_ & new_n_n31_;
  assign new_nmis15847_ = new_nmis16866_ & new_nxz324_ & new_nmis11550_ & new_nenwin_ & new_nmis16858_ & new_nmis16864_;
  assign new_n_n117_ = new_nmis16657_ & new_nslad0_;
  assign new_nmis16889_ = new_nvzzze_ | new_n_n44_;
  assign new_nmis11562_ = new_n_n47_ & new_nvfin_;
  assign new_nmis16716_ = new_n_n91_ | new_n_n92_;
  assign new_n_n87_ = new_naxz1_ & new_n_n55_;
  assign new_n_n2_ = ~new_nmis16883_;
  assign new_n_n382_ = new_nxzfr1_ & new_n_n22_;
  assign new_np1zzz3_p_ = new_n_n373_ | new_n_n374_;
  assign new_n_n352_ = new_nmis11585_ & new_np2zzz6_;
  assign new_ni1zzz2_p_ = new_n_n343_ | new_n_n344_;
  assign new_n_n340_ = new_nmis11581_ & new_ni1zzz4_;
  assign new_ni2zzz0_p_ = new_n_n331_ | new_n_n332_;
  assign new_n_n328_ = new_nmis11583_ & new_ni2zzz2_;
  assign new_ni2zzz6_p_ = new_n_n319_ | new_n_n320_;
  assign new_nryz_p_ = new_n_n221_ | new_niclr_;
  assign new_n_n312_ = new_nmis8641_ & new_n_n32_;
  assign new_nqpr2_p_ = new_n_n303_ | new_n_n304_;
  assign new_n_n294_ = new_nmis11589_ & new_nv1zzz2_;
  assign new_nv1zzz6_p_ = new_n_n285_ | new_n_n286_;
  assign new_n_n282_ = new_nmis11591_ & new_nv2zzz0_;
  assign new_nv2zzz4_p_ = new_n_n273_ | new_n_n274_;
  assign new_n_n270_ = new_nmis11591_ & new_nv2zzz6_;
  assign new_n_n263_ = new_ni1zzz2_ & new_nmis11594_;
  assign new_n_n258_ = new_np1zzz4_ & new_nmis15081_;
  assign new_ntxwrd8_p_ = new_n_n250_ | new_n_n249_ | new_n_n248_;
  assign new_n_n241_ = new_ni2zzz6_ & new_nmis11594_;
  assign new_n_n234_ = new_nxz321_ & new_n_n50_ & new_nmis15083_;
  assign new_nxz160_f_ = new_n_n228_ | new_n_n229_;
  assign new_n_n222_ = new_nmis15848_ & new_n_n63_ & new_nmis11560_ & new_nxz162_;
  assign new_n_n219_ = new_nrptwin_ & new_nrpten_ & new_nmis16712_;
  assign new_nmis11556_ = new_n_n30_ & new_naxz0_ & new_naxz1_;
  assign new_n_n213_ = new_n_n68_ & new_n_n70_ & new_n_n6_;
  assign new_n_n209_ = new_n_n22_ & new_nmis16752_;
  assign new_nmis16748_ = new_n_n204_ | new_na_;
  assign new_nmis16548_ = new_nmis16581_ | new_n_n41_;
  assign new_nmis11593_ = new_n_n19_ & new_n_n46_;
  assign new_n_n185_ = new_nmis11562_ & new_nv1zzz2_;
  assign new_nmis16728_ = new_n_n181_ | new_n_n180_ | new_n_n179_;
  assign new_n_n173_ = new_nmis11549_ & new_ntxwrd7_;
  assign new_n_n168_ = new_nmis11548_ & new_ntxwrd8_;
  assign new_nmis16596_ = new_n_n159_ | new_n_n158_ | new_n_n157_;
  assign new_n_n154_ = new_ni2zzz4_ & new_ninfin_;
  assign new_n_n146_ = new_nmis15062_ & new_ntxwrd15_;
  assign new_n_n139_ = new_nmis11560_ & new_n_n56_;
  assign new_n_n129_ = new_n_n55_ & new_nrxz0_ & new_n_n33_;
  assign new_nmis16572_ = new_n_n124_ | new_ntxmess_n_;
  assign new_nmis7564_ = new_n_n51_ | new_n_n34_ | new_n_n35_;
  assign new_nmis15328_ = new_n_n115_ | new_n_n71_;
  assign new_nmis9061_ = new_n_n112_ | new_ntxmess_n_;
  assign new_nmis15065_ = new_nmis11549_ & new_n_n47_;
  assign new_n_n106_ = new_nmis11549_ & new_ntxwrd8_;
  assign new_n_n98_ = new_nmis11548_ & new_ntxwrd12_;
  assign new_n_n3_ = ~new_nmis16885_;
  assign new_n_n381_ = new_nofs2_p_ & new_nofs2_;
  assign new_n_n375_ = new_nmis11588_ & new_npybb3_;
  assign new_n_n351_ = new_nmis11586_ & new_npybb7_;
  assign new_n_n345_ = new_nmis11582_ & new_ninybb2_;
  assign new_n_n339_ = new_nmis11582_ & new_ninybb5_;
  assign new_n_n333_ = new_nmis11582_ & new_ninybb8_;
  assign new_n_n327_ = new_nmis11584_ & new_ninybb3_;
  assign new_n_n321_ = new_nmis11584_ & new_ninybb6_;
  assign new_ncomppar_p_ = new_n_n19_ & new_nmis16569_;
  assign new_nrxz0_p_ = new_n_n311_ | new_n_n312_;
  assign new_naxz1_p_ = new_n_n19_ & new_nmis16553_;
  assign new_n_n293_ = new_nmis11590_ & new_nv1zzz3_;
  assign new_n_n287_ = new_nmis11590_ & new_nv1zzz6_;
  assign new_n_n281_ = new_nmis11592_ & new_nv2zzz1_;
  assign new_n_n275_ = new_nmis11592_ & new_nv2zzz4_;
  assign new_n_n269_ = new_nmis11592_ & new_nv2zzz7_;
  assign new_n_n264_ = new_nmis16585_ & new_nmis11593_;
  assign new_n_n257_ = new_nmis15080_ & new_nmis16728_;
  assign new_ntxwrd7_p_ = new_n_n19_ & new_nmis16618_;
  assign new_n_n240_ = new_nmis15080_ & new_nmis16736_;
  assign new_n_n235_ = new_nmis15339_ & new_nxz322_;
  assign new_n_n229_ = new_nmis16754_ & new_nxz160_n_;
  assign new_n_n223_ = new_nmis16602_ & new_nxz163_;
  assign new_n_n218_ = new_nmis16690_ & new_n_n42_ & new_nmis16710_ & new_n_n58_;
  assign new_nmis11565_ = new_ntxmess_n_ & new_n_n49_ & new_nmis11547_;
  assign new_nmis10130_ = new_n_n212_ | new_nxz320_p_;
  assign new_nmis8641_ = new_n_n208_ | new_n_n209_;
  assign new_n_n204_ = new_n_n10_ & new_n_n30_;
  assign new_nmis15843_ = new_nqpr1_ & new_nqpr0_ & new_n_n15_;
  assign new_nmis11594_ = new_n_n19_ & new_ninfin_;
  assign new_n_n186_ = new_nmis15065_ & new_ntxwrd3_;
  assign new_n_n181_ = new_nv1zzz4_ & new_nvfin_;
  assign new_n_n174_ = new_nmis11548_ & new_ntxwrd6_;
  assign new_n_n167_ = new_nmis11549_ & new_ntxwrd9_;
  assign new_n_n160_ = new_ni2zzz2_ & new_ninfin_;
  assign new_nmis16734_ = new_n_n153_ | new_n_n152_ | new_n_n151_;
  assign new_n_n147_ = new_np2zzz7_ & new_npfin_;
  assign new_nmis11550_ = new_nxz320_ & new_nxz323_ & new_nmis11578_;
  assign new_nmis16883_ = new_npzzze_ | new_n_n26_;
  assign new_n_n125_ = new_nmis16577_ & new_n_n30_ & new_n_n62_;
  assign new_nmis16752_ = new_nmis15847_ | new_nrptwin_;
  assign new_nmis16765_ = new_n_n38_ | new_nmis8768_;
  assign new_n_n112_ = new_nmis16765_ & new_n_n43_;
  assign new_nmis15062_ = new_nmis11548_ & new_n_n47_;
  assign new_nmis16611_ = new_n_n105_ | new_n_n104_ | new_n_n103_;
  assign new_n_n99_ = new_nv2zzz4_ & new_nvfin_;
  assign new_n_n4_ = ~new_nmis16891_;
  assign new_nmis16746_ = new_n_n81_ | new_n_n82_;
  assign new_nmis16873_ = new_n_n75_ | new_n_n76_;
  assign new_n_n72_ = ~new_nb_;
  assign new_n_n61_ = ~new_naxz0_;
  assign new_n_n50_ = ~new_nxz322_;
  assign new_nmis12425_ = new_nmis16673_ | new_n_n57_;
  assign new_n_n76_ = new_nslad2_ & new_nxz162_;
  assign new_nmis16767_ = new_n_n72_ | new_nqpr4_;
  assign new_n_n60_ = ~new_nmis9255_;
  assign new_n_n51_ = ~new_nxz323_;
  assign new_nmis16657_ = new_nmis10125_ | new_nmis16027_ | new_nmis12425_;
  assign new_n_n75_ = new_n_n65_ & new_n_n64_;
  assign new_n_n70_ = ~new_nslad1_;
  assign new_n_n63_ = ~new_nxz163_;
  assign new_n_n52_ = ~new_nqpr0_;
  assign new_nmis16675_ = new_nmis16027_ | new_nmis16023_;
  assign new_nmis15855_ = new_nxz162_ & new_n_n65_;
  assign new_n_n71_ = ~new_ncbt2_;
  assign new_n_n62_ = ~new_ncomppar_;
  assign new_n_n53_ = ~new_naxz1_;
  assign new_n_n0_ = ~new_nmis8027_;
  assign new_nmis16673_ = new_nmis15855_ | new_nmis15854_;
  assign new_n_n43_ = ~new_na_;
  assign new_n_n32_ = ~new_nrxz0_;
  assign new_n_n21_ = ~new_nmis10125_;
  assign new_n_n10_ = ~new_nmis16765_;
  assign new_nmis16646_ = new_n_n69_ | new_nmis12425_ | new_n_n56_ | new_nmis16023_;
  assign new_n_n42_ = ~new_nqpr4_;
  assign new_n_n33_ = ~new_nrxz1_;
  assign new_n_n20_ = ~new_nxz321_;
  assign new_n_n11_ = ~new_nmis8768_;
  assign new_n_n41_ = ~new_nqpr2_;
  assign new_n_n30_ = ~new_ntxmess_n_;
  assign new_n_n23_ = ~new_nqpr1_;
  assign new_n_n12_ = ~new_nmis15328_;
  assign new_n_n40_ = ~new_ncbt0_;
  assign new_n_n31_ = ~new_nmis11154_;
  assign new_n_n22_ = ~new_niclr_;
  assign new_n_n13_ = ~new_nmis9174_;
  assign new_n_n69_ = ~new_nenwin_;
  assign new_n_n58_ = ~new_nqpr3_;
  assign new_n_n47_ = ~new_npfin_;
  assign new_n_n36_ = ~new_npsync_;
  assign new_n_n25_ = ~new_nrptwin_;
  assign new_n_n14_ = ~new_nc_;
  assign new_n_n68_ = ~new_nslad0_;
  assign new_n_n59_ = ~new_nmis16767_;
  assign new_n_n46_ = ~new_ninfin_;
  assign new_n_n37_ = ~new_nxzfs_;
  assign new_n_n24_ = ~new_nsbuff_;
  assign new_n_n15_ = ~new_ntxmess_f_;
  assign new_nmis16719_ = new_n_n79_ | new_n_n80_;
  assign new_nmis16023_ = new_n_n74_ | new_nmis7564_;
  assign new_n_n45_ = ~new_nvzzze_;
  assign new_n_n34_ = ~new_nxz324_;
  assign new_n_n27_ = ~new_npzzze_;
  assign new_n_n16_ = ~new_nmis9061_;
  assign new_n_n80_ = new_n_n61_ & new_nesrsum_;
  assign new_nmis15854_ = new_nxz163_ & new_n_n66_;
  assign new_n_n44_ = ~new_nvybb0_;
  assign new_n_n35_ = ~new_nmis11578_;
  assign new_n_n26_ = ~new_npybb0_;
  assign new_n_n17_ = ~new_nmis16889_;
  assign new_nmis16792_ = new_n_n60_ | new_ntxmess_n_;
  assign new_n_n79_ = new_n_n62_ & new_naxz0_;
  assign new_nmis16027_ = new_n_n73_ | new_n_n69_;
  assign new_n_n65_ = ~new_nslad2_;
  assign new_n_n54_ = ~new_nmmerr_;
  assign new_n_n29_ = ~new_ninzzze_;
  assign new_n_n18_ = ~new_nmis16893_;
  assign new_nmis16895_ = new_ncbt0_ | new_ncbt1_ | new_n_n71_;
  assign new_nmis16871_ = new_n_n77_ | new_n_n78_;
  assign new_n_n74_ = new_n_n67_ & new_n_n68_;
  assign new_n_n64_ = ~new_nxz162_;
  assign new_n_n55_ = ~new_nesrsum_;
  assign new_n_n28_ = ~new_ninybb0_;
  assign new_n_n19_ = ~new_nryz_;
  assign new_n_n81_ = new_n_n59_ & new_nqpr3_;
  assign new_n_n78_ = new_nxz163_ & new_nslad3_;
  assign new_nmis16750_ = new_nqpr4_ | new_n_n71_;
  assign new_n_n67_ = ~new_nxz160_n_;
  assign new_n_n56_ = ~new_nxz161_;
  assign new_n_n49_ = ~new_nvfin_;
  assign new_n_n38_ = ~new_nmis16746_;
  assign new_n_n82_ = new_n_n58_ & new_nmis16750_;
  assign new_n_n77_ = new_n_n63_ & new_n_n66_;
  assign new_n_n73_ = new_nxz161_ & new_n_n70_;
  assign new_n_n66_ = ~new_nslad3_;
  assign new_n_n57_ = ~new_nxz320_;
  assign new_n_n48_ = ~new_nmis16792_;
  assign new_n_n39_ = ~new_ncbt1_;
endmodule


