// Benchmark "top" written by ABC on Fri Mar 31 12:09:39 2023

module top ( 
    pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps, pd0, pe1,
    pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0, pw, ph0,
    pi1, px, ph1, pi0, py, ph2, pj0, pk1, pz, pj1, pk0, pl0, pm1, pl1, pm0,
    pn0, po1, pn1, po0, pp0, pq1, pa, pp1, pq0, pb, pr0, ps1, pr1, ps0, pd,
    pt0, pu1, pe, pt1, pu0, pf, pv0, pw1, pg, pv1, pw0, ph, px0, py1, pi,
    px1, py0, pj, pz0, pk, pz1, pl, pm, pn, po,
    pc3, pd4, pb3, pe4, pa3, pf4, pg4, pg3, pa4, pf3, pb4, pe3, pc4, pd3,
    pj2, pk3, pl4, pj3, pk2, pm4, pi3, pn4, ph3, pi2, po4, ph4, pn2, po3,
    pi4, pn3, po2, pj4, pl2, pm3, pk4, pl3, pm2, pr2, ps3, pt4, pr3, ps2,
    pu4, pp2, pq3, pv4, pp3, pq2, pp4, pv2, pw3, pq4, pv3, pw2, pr4, pt2,
    pu3, ps4, pt3, pu2, pz2, pz3, px2, py3, px3, py2  );
  input  pa1, pb2, pp, pa0, pc2, pq, pb0, pc1, pr, pa2, pb1, pc0, ps,
    pd0, pe1, pf2, pt, pd1, pe0, pg2, pu, pd2, pf0, pg1, pv, pe2, pf1, pg0,
    pw, ph0, pi1, px, ph1, pi0, py, ph2, pj0, pk1, pz, pj1, pk0, pl0, pm1,
    pl1, pm0, pn0, po1, pn1, po0, pp0, pq1, pa, pp1, pq0, pb, pr0, ps1,
    pr1, ps0, pd, pt0, pu1, pe, pt1, pu0, pf, pv0, pw1, pg, pv1, pw0, ph,
    px0, py1, pi, px1, py0, pj, pz0, pk, pz1, pl, pm, pn, po;
  output pc3, pd4, pb3, pe4, pa3, pf4, pg4, pg3, pa4, pf3, pb4, pe3, pc4, pd3,
    pj2, pk3, pl4, pj3, pk2, pm4, pi3, pn4, ph3, pi2, po4, ph4, pn2, po3,
    pi4, pn3, po2, pj4, pl2, pm3, pk4, pl3, pm2, pr2, ps3, pt4, pr3, ps2,
    pu4, pp2, pq3, pv4, pp3, pq2, pp4, pv2, pw3, pq4, pv3, pw2, pr4, pt2,
    pu3, ps4, pt3, pu2, pz2, pz3, px2, py3, px3, py2;
  wire new_na1_, new_nb2_, new_np_, new_na0_, new_nc2_, new_nq_, new_nb0_,
    new_nc1_, new_nr_, new_na2_, new_nb1_, new_nc0_, new_ns_, new_nd0_,
    new_ne1_, new_nf2_, new_nt_, new_nd1_, new_ne0_, new_ng2_, new_nu_,
    new_nd2_, new_nf0_, new_ng1_, new_nv_, new_ne2_, new_nf1_, new_ng0_,
    new_nw_, new_nh0_, new_ni1_, new_nx_, new_nh1_, new_ni0_, new_ny_,
    new_nh2_, new_nj0_, new_nk1_, new_nz_, new_nj1_, new_nk0_, new_nl0_,
    new_nm1_, new_nl1_, new_nm0_, new_nn0_, new_no1_, new_nn1_, new_no0_,
    new_np0_, new_nq1_, new_na_, new_np1_, new_nq0_, new_nb_, new_nr0_,
    new_ns1_, new_nr1_, new_ns0_, new_nd_, new_nt0_, new_nu1_, new_ne_,
    new_nt1_, new_nu0_, new_nf_, new_nv0_, new_nw1_, new_ng_, new_nv1_,
    new_nw0_, new_nh_, new_nx0_, new_ny1_, new_ni_, new_nx1_, new_ny0_,
    new_nj_, new_nz0_, new_nk_, new_nz1_, new_nl_, new_nm_, new_nn_,
    new_no_, new_n_n137_, new_n_n131_, new_ns2_, new_ni3_, new_nr3_,
    new_nc4_, new_n_n85_, new_n_n77_, new_n_n69_, new_n_n138_, new_n_n130_,
    new_n_n124_, new_nj3_, new_nq3_, new_nd4_, new_n_n86_, new_n_n76_,
    new_nk4_, new_n_n136_, new_n_n132_, new_n_n125_, new_na3_, new_n_n100_,
    new_n_n93_, new_n_n84_, new_nh4_, new_n_n70_, new_nk2_, new_no2_,
    new_nr2_, new_n_n107_, new_n_n101_, new_n_n92_, new_nf4_, new_n_n78_,
    new_n_n71_, new_ni2_, new_nl2_, new_n_n128_, new_n_n121_, new_nx2_,
    new_n_n91_, new_n_n82_, new_n_n74_, new_n_n67_, new_n_n9_, new_n_n142_,
    new_n_n135_, new_nt2_, new_n_n120_, new_n_n114_, new_n_n90_,
    new_n_n83_, new_n_n73_, new_nm4_, new_n_n141_, new_np2_, new_n_n122_,
    new_n_n89_, new_n_n81_, new_ni4_, new_nl4_, new_nm2_, new_n_n129_,
    new_n_n123_, new_n_n88_, new_ng4_, new_n_n75_, new_n_n68_, new_n_n118_,
    new_n_n111_, new_nc3_, new_n_n97_, new_n_n95_, new_nz3_, new_n_n5_,
    new_nv2_, new_ny2_, new_n_n103_, new_ng3_, new_n_n94_, new_ny3_,
    new_n_n6_, new_nu2_, new_n_n112_, new_n_n102_, new_nh3_, new_no3_,
    new_nx3_, new_n_n7_, new_n_n119_, new_n_n113_, new_nd3_, new_n_n96_,
    new_np3_, new_nw3_, new_n_n8_, new_n_n140_, new_nn2_, new_n_n126_,
    new_nw2_, new_n_n108_, new_n_n106_, new_n_n99_, new_nm3_, new_nv3_,
    new_n_n80_, new_n_n72_, new_n_n1_, new_n_n133_, new_n_n127_,
    new_n_n115_, new_n_n109_, new_nb3_, new_ne3_, new_nn3_, new_nu3_,
    new_n_n79_, new_nj4_, new_n_n2_, new_n_n139_, new_nq2_, new_n_n117_,
    new_nz2_, new_n_n105_, new_n_n98_, new_nk3_, new_nt3_, new_na4_,
    new_n_n87_, new_n_n3_, new_nj2_, new_n_n134_, new_n_n116_, new_n_n110_,
    new_n_n104_, new_nf3_, new_nl3_, new_ns3_, new_nb4_, new_ne4_,
    new_n_n4_, new_nn4_, new_nq4_, new_ns4_, new_n_n39_, new_ng10_,
    new_n_n62_, new_n_n53_, new_n_n45_, new_na10_, new_nf10_, new_n_n63_,
    new_n_n52_, new_nt4_, new_nz9_, new_ne10_, new_n_n64_, new_n_n51_,
    new_n_n44_, new_n_n40_, new_n_n35_, new_n_n0_, new_n_n65_, new_n_n30_,
    new_nr10_, new_n_n21_, new_n_n10_, new_n_n66_, new_nj10_, new_nq10_,
    new_n_n20_, new_n_n11_, new_nk10_, new_ns10_, new_n_n23_, new_n_n12_,
    new_nl10_, new_n_n27_, new_n_n22_, new_n_n13_, new_nu4_, new_n_n38_,
    new_nh10_, new_nn10_, new_nv10_, new_n_n14_, new_n_n43_, new_nb10_,
    new_ni10_, new_n_n28_, new_n_n24_, new_n_n15_, new_n_n58_, new_n_n49_,
    new_n_n32_, new_np10_, new_nt10_, new_n_n16_, new_n_n57_, new_n_n50_,
    new_n_n31_, new_no10_, new_nu10_, new_n_n17_, new_n_n59_, new_np4_,
    new_nr4_, new_ny9_, new_n_n36_, new_n_n26_, new_n_n18_, new_n_n60_,
    new_n_n56_, new_n_n48_, new_n_n41_, new_nd10_, new_n_n25_, new_n_n19_,
    new_n_n61_, new_n_n55_, new_n_n46_, new_n_n42_, new_nc10_, new_n_n34_,
    new_n_n29_, new_no4_, new_n_n54_, new_n_n47_, new_nv4_, new_n_n37_,
    new_n_n33_, new_nm10_;
  assign new_na1_ = pa1;
  assign new_nb2_ = pb2;
  assign pc3 = new_nc3_;
  assign pd4 = new_nd4_;
  assign new_np_ = pp;
  assign new_na0_ = pa0;
  assign pb3 = new_nb3_;
  assign new_nc2_ = pc2;
  assign pe4 = new_ne4_;
  assign new_nq_ = pq;
  assign pa3 = new_na3_;
  assign new_nb0_ = pb0;
  assign new_nc1_ = pc1;
  assign pf4 = new_nf4_;
  assign new_nr_ = pr;
  assign new_na2_ = pa2;
  assign new_nb1_ = pb1;
  assign new_nc0_ = pc0;
  assign pg4 = new_ng4_;
  assign new_ns_ = ps;
  assign new_nd0_ = pd0;
  assign new_ne1_ = pe1;
  assign new_nf2_ = pf2;
  assign pg3 = new_ng3_;
  assign new_nt_ = pt;
  assign pa4 = new_na4_;
  assign new_nd1_ = pd1;
  assign new_ne0_ = pe0;
  assign pf3 = new_nf3_;
  assign new_ng2_ = pg2;
  assign new_nu_ = pu;
  assign pb4 = new_nb4_;
  assign new_nd2_ = pd2;
  assign pe3 = new_ne3_;
  assign new_nf0_ = pf0;
  assign new_ng1_ = pg1;
  assign new_nv_ = pv;
  assign pc4 = new_nc4_;
  assign pd3 = new_nd3_;
  assign new_ne2_ = pe2;
  assign new_nf1_ = pf1;
  assign new_ng0_ = pg0;
  assign new_nw_ = pw;
  assign new_nh0_ = ph0;
  assign new_ni1_ = pi1;
  assign pj2 = new_nj2_;
  assign pk3 = new_nk3_;
  assign pl4 = new_nl4_;
  assign new_nx_ = px;
  assign new_nh1_ = ph1;
  assign new_ni0_ = pi0;
  assign pj3 = new_nj3_;
  assign pk2 = new_nk2_;
  assign pm4 = new_nm4_;
  assign new_ny_ = py;
  assign new_nh2_ = ph2;
  assign pi3 = new_ni3_;
  assign new_nj0_ = pj0;
  assign new_nk1_ = pk1;
  assign pn4 = new_nn4_;
  assign new_nz_ = pz;
  assign ph3 = new_nh3_;
  assign pi2 = new_ni2_;
  assign new_nj1_ = pj1;
  assign new_nk0_ = pk0;
  assign po4 = new_no4_;
  assign ph4 = new_nh4_;
  assign new_nl0_ = pl0;
  assign new_nm1_ = pm1;
  assign pn2 = new_nn2_;
  assign po3 = new_no3_;
  assign pi4 = new_ni4_;
  assign new_nl1_ = pl1;
  assign new_nm0_ = pm0;
  assign pn3 = new_nn3_;
  assign po2 = new_no2_;
  assign pj4 = new_nj4_;
  assign pl2 = new_nl2_;
  assign pm3 = new_nm3_;
  assign new_nn0_ = pn0;
  assign new_no1_ = po1;
  assign pk4 = new_nk4_;
  assign pl3 = new_nl3_;
  assign pm2 = new_nm2_;
  assign new_nn1_ = pn1;
  assign new_no0_ = po0;
  assign new_np0_ = pp0;
  assign new_nq1_ = pq1;
  assign pr2 = new_nr2_;
  assign ps3 = new_ns3_;
  assign pt4 = new_nt4_;
  assign new_na_ = pa;
  assign new_np1_ = pp1;
  assign new_nq0_ = pq0;
  assign pr3 = new_nr3_;
  assign ps2 = new_ns2_;
  assign pu4 = new_nu4_;
  assign new_nb_ = pb;
  assign pp2 = new_np2_;
  assign pq3 = new_nq3_;
  assign new_nr0_ = pr0;
  assign new_ns1_ = ps1;
  assign pv4 = new_nv4_;
  assign pp3 = new_np3_;
  assign pq2 = new_nq2_;
  assign new_nr1_ = pr1;
  assign new_ns0_ = ps0;
  assign new_nd_ = pd;
  assign pp4 = new_np4_;
  assign new_nt0_ = pt0;
  assign new_nu1_ = pu1;
  assign pv2 = new_nv2_;
  assign pw3 = new_nw3_;
  assign new_ne_ = pe;
  assign pq4 = new_nq4_;
  assign new_nt1_ = pt1;
  assign new_nu0_ = pu0;
  assign pv3 = new_nv3_;
  assign pw2 = new_nw2_;
  assign new_nf_ = pf;
  assign pr4 = new_nr4_;
  assign pt2 = new_nt2_;
  assign pu3 = new_nu3_;
  assign new_nv0_ = pv0;
  assign new_nw1_ = pw1;
  assign new_ng_ = pg;
  assign ps4 = new_ns4_;
  assign pt3 = new_nt3_;
  assign pu2 = new_nu2_;
  assign new_nv1_ = pv1;
  assign new_nw0_ = pw0;
  assign new_nh_ = ph;
  assign new_nx0_ = px0;
  assign new_ny1_ = py1;
  assign pz2 = new_nz2_;
  assign new_ni_ = pi;
  assign new_nx1_ = px1;
  assign new_ny0_ = py0;
  assign pz3 = new_nz3_;
  assign new_nj_ = pj;
  assign px2 = new_nx2_;
  assign py3 = new_ny3_;
  assign new_nz0_ = pz0;
  assign new_nk_ = pk;
  assign px3 = new_nx3_;
  assign py2 = new_ny2_;
  assign new_nz1_ = pz1;
  assign new_nl_ = pl;
  assign new_nm_ = pm;
  assign new_nn_ = pn;
  assign new_no_ = po;
  assign new_n_n137_ = new_n_n15_ & new_n_n13_ & new_n_n10_;
  assign new_n_n131_ = new_n_n5_ & new_nz_;
  assign new_ns2_ = new_n_n122_ | new_n_n123_;
  assign new_ni3_ = new_nz9_ & new_nt0_;
  assign new_nr3_ = new_ny9_ & new_nc1_;
  assign new_nc4_ = new_ny9_ & new_nn1_;
  assign new_n_n85_ = new_nq10_ & new_nr1_;
  assign new_n_n77_ = new_np10_ & new_nm_;
  assign new_n_n69_ = new_no10_ & new_nx_;
  assign new_n_n138_ = new_n_n9_ & new_n_n15_;
  assign new_n_n130_ = new_nn1_ & new_np0_;
  assign new_n_n124_ = new_nk1_ & new_np0_;
  assign new_nj3_ = new_nz9_ & new_nu0_;
  assign new_nq3_ = new_ny9_ & new_nb1_;
  assign new_nd4_ = new_n_n88_ | new_n_n91_ | new_n_n93_ | new_n_n92_ | new_n_n90_ | new_n_n89_;
  assign new_n_n86_ = new_np10_ & new_nj_;
  assign new_n_n76_ = new_nq10_ & new_nu1_;
  assign new_nk4_ = new_n_n68_ | new_n_n69_;
  assign new_n_n136_ = new_nh10_ & new_np1_ & new_nj10_;
  assign new_n_n132_ = new_no1_ & new_np0_;
  assign new_n_n125_ = new_n_n5_ & new_nc0_;
  assign new_na3_ = new_n_n106_ | new_n_n107_;
  assign new_n_n100_ = new_nt0_ & new_np0_;
  assign new_n_n93_ = new_ni_ & new_np10_;
  assign new_n_n84_ = new_no10_ & new_ns_;
  assign new_nh4_ = new_n_n78_ | new_n_n77_ | new_n_n76_;
  assign new_n_n70_ = new_nq10_ & new_nw1_;
  assign new_nk2_ = new_n_n135_ | new_n_n136_;
  assign new_no2_ = new_n_n130_ | new_n_n131_;
  assign new_nr2_ = new_n_n124_ | new_n_n125_;
  assign new_n_n107_ = new_n_n5_ & new_nl0_;
  assign new_n_n101_ = new_n_n5_ & new_no0_;
  assign new_n_n92_ = new_nq_ & new_no10_;
  assign new_nf4_ = new_n_n84_ | new_n_n83_ | new_n_n82_;
  assign new_n_n78_ = new_no10_ & new_nu_;
  assign new_n_n71_ = new_np10_ & new_no_;
  assign new_ni2_ = new_n_n142_ | new_n_n141_ | new_n_n140_;
  assign new_nl2_ = new_nb1_ & new_n_n15_ & new_nl10_;
  assign new_n_n128_ = new_nm1_ & new_np0_;
  assign new_n_n121_ = new_n_n5_ & new_ne0_;
  assign new_nx2_ = new_n_n112_ | new_n_n113_;
  assign new_n_n91_ = new_nj10_ & new_nc2_ & new_n_n15_ & new_n_n16_ & new_nq1_;
  assign new_n_n82_ = new_nq10_ & new_ns1_;
  assign new_n_n74_ = new_np10_ & new_nn_;
  assign new_n_n67_ = new_n_n10_ & new_n_n13_;
  assign new_n_n9_ = ~new_nc10_;
  assign new_n_n142_ = new_n_n5_ & new_nh_;
  assign new_n_n135_ = new_nh10_ & new_ny1_ & new_nk10_;
  assign new_nt2_ = new_n_n120_ | new_n_n121_;
  assign new_n_n120_ = new_ni1_ & new_np0_;
  assign new_n_n114_ = new_na1_ & new_np0_;
  assign new_n_n90_ = new_nj10_ & new_nc2_ & new_n_n15_ & new_n_n16_ & new_ny1_;
  assign new_n_n83_ = new_np10_ & new_nk_;
  assign new_n_n73_ = new_nq10_ & new_nv1_;
  assign new_nm4_ = new_n_n64_ | new_n_n63_ | new_nb_ | new_n_n62_ | new_n_n66_ | new_n_n65_ | new_n_n1_ | new_n_n67_;
  assign new_n_n141_ = new_nb1_ & new_np0_;
  assign new_np2_ = new_n_n128_ | new_n_n129_;
  assign new_n_n122_ = new_nj1_ & new_np0_;
  assign new_n_n89_ = new_nq0_ & new_nd2_ & new_np1_ & new_nj10_ & new_nc2_ & new_n_n15_ & new_ne10_ & new_nd10_;
  assign new_n_n81_ = new_no10_ & new_nt_;
  assign new_ni4_ = new_n_n75_ | new_n_n74_ | new_n_n73_;
  assign new_nl4_ = new_n_n21_ & new_nh2_ & new_ng2_ & new_na10_ & new_nv10_;
  assign new_nm2_ = new_n_n134_ | new_nh10_;
  assign new_n_n129_ = new_n_n5_ & new_na0_;
  assign new_n_n123_ = new_n_n5_ & new_nd0_;
  assign new_n_n88_ = new_n_n3_ & new_nd2_ & new_n_n0_ & new_nj10_ & new_nc2_ & new_n_n15_ & new_ne10_ & new_nd10_;
  assign new_ng4_ = new_n_n81_ | new_n_n80_ | new_n_n79_;
  assign new_n_n75_ = new_no10_ & new_nv_;
  assign new_n_n68_ = new_np10_ & new_np_;
  assign new_n_n118_ = new_nh1_ & new_np0_;
  assign new_n_n111_ = new_n_n5_ & new_nj0_;
  assign new_nc3_ = new_n_n102_ | new_n_n103_;
  assign new_n_n97_ = new_n_n15_ & new_n_n12_ & new_ng_ & new_n_n20_ & new_n_n11_;
  assign new_n_n95_ = new_nz9_ & new_na1_;
  assign new_nz3_ = new_ny9_ & new_nk1_;
  assign new_n_n5_ = ~new_np0_;
  assign new_nv2_ = new_n_n116_ | new_n_n117_;
  assign new_ny2_ = new_n_n110_ | new_n_n111_;
  assign new_n_n103_ = new_n_n5_ & new_nn0_;
  assign new_ng3_ = new_n_n96_ | new_n_n97_;
  assign new_n_n94_ = new_ng_ & new_nb10_ & new_nr0_ & new_na10_;
  assign new_ny3_ = new_ny9_ & new_nj1_;
  assign new_n_n6_ = ~new_nu10_;
  assign new_nu2_ = new_n_n118_ | new_n_n119_;
  assign new_n_n112_ = new_nz0_ & new_np0_;
  assign new_n_n102_ = new_nu0_ & new_np0_;
  assign new_nh3_ = new_nz9_ & new_ng_;
  assign new_no3_ = new_nz9_ & new_nz0_;
  assign new_nx3_ = new_ny9_ & new_ni1_;
  assign new_n_n7_ = ~new_ne10_;
  assign new_n_n119_ = new_n_n5_ & new_nf0_;
  assign new_n_n113_ = new_n_n5_ & new_ni0_;
  assign new_nd3_ = new_n_n100_ | new_n_n101_;
  assign new_n_n96_ = new_n_n15_ & new_n_n12_ & new_ng_ & new_n_n20_ & new_n_n9_;
  assign new_np3_ = new_n_n94_ | new_n_n95_;
  assign new_nw3_ = new_ny9_ & new_nh1_;
  assign new_n_n8_ = ~new_ns10_;
  assign new_n_n140_ = new_nm2_ & new_np0_;
  assign new_nn2_ = new_n_n132_ | new_n_n133_;
  assign new_n_n126_ = new_nl1_ & new_np0_;
  assign new_nw2_ = new_n_n114_ | new_n_n115_;
  assign new_n_n108_ = new_nx0_ & new_np0_;
  assign new_n_n106_ = new_nw0_ & new_np0_;
  assign new_n_n99_ = new_n_n3_ & new_nk2_ & new_n_n16_;
  assign new_nm3_ = new_nz9_ & new_nx0_;
  assign new_nv3_ = new_ny9_ & new_ng1_;
  assign new_n_n80_ = new_np10_ & new_nl_;
  assign new_n_n72_ = new_no10_ & new_nw_;
  assign new_n_n1_ = ~new_na_;
  assign new_n_n133_ = new_n_n5_ & new_ny_;
  assign new_n_n127_ = new_n_n5_ & new_nb0_;
  assign new_n_n115_ = new_n_n5_ & new_nh0_;
  assign new_n_n109_ = new_n_n5_ & new_nk0_;
  assign new_nb3_ = new_n_n104_ | new_n_n105_;
  assign new_ne3_ = new_n_n99_ | new_ng10_;
  assign new_nn3_ = new_nz9_ & new_ny0_;
  assign new_nu3_ = new_ny9_ & new_nf1_;
  assign new_n_n79_ = new_nq10_ & new_nt1_;
  assign new_nj4_ = new_n_n72_ | new_n_n71_ | new_n_n70_;
  assign new_n_n2_ = ~new_ny1_;
  assign new_n_n139_ = new_n_n11_ & new_n_n15_;
  assign new_nq2_ = new_n_n126_ | new_n_n127_;
  assign new_n_n117_ = new_n_n5_ & new_ng0_;
  assign new_nz2_ = new_n_n108_ | new_n_n109_;
  assign new_n_n105_ = new_n_n5_ & new_nm0_;
  assign new_n_n98_ = new_ng_ & new_n_n12_ & new_n_n11_;
  assign new_nk3_ = new_nz9_ & new_nv0_;
  assign new_nt3_ = new_ny9_ & new_ne1_;
  assign new_na4_ = new_ny9_ & new_nl1_;
  assign new_n_n87_ = new_no10_ & new_nr_;
  assign new_n_n3_ = ~new_nq0_;
  assign new_nj2_ = new_n_n139_ | new_n_n138_ | new_n_n137_;
  assign new_n_n134_ = new_nc10_ & new_n_n15_;
  assign new_n_n116_ = new_ng1_ & new_np0_;
  assign new_n_n110_ = new_ny0_ & new_np0_;
  assign new_n_n104_ = new_nv0_ & new_np0_;
  assign new_nf3_ = new_n_n1_ | new_nb_ | new_n_n98_;
  assign new_nl3_ = new_nz9_ & new_nw0_;
  assign new_ns3_ = new_ny9_ & new_nd1_;
  assign new_nb4_ = new_ny9_ & new_nm1_;
  assign new_ne4_ = new_n_n87_ | new_n_n86_ | new_n_n85_;
  assign new_n_n4_ = ~new_nd_;
  assign new_nn4_ = new_na_ & new_n_n4_ & new_ne_ & new_n_n15_;
  assign new_nq4_ = new_n_n48_ | new_n_n51_ | new_n_n53_ | new_n_n52_ | new_n_n50_ | new_n_n49_;
  assign new_ns4_ = new_n_n44_ | new_ng10_;
  assign new_n_n39_ = new_na10_ & new_n_n22_ & new_n_n17_ & new_n_n19_;
  assign new_ng10_ = new_n_n33_ | new_n_n34_;
  assign new_n_n62_ = new_n_n13_ & new_nd10_ & new_nc2_ & new_n_n3_ & new_n_n2_;
  assign new_n_n53_ = new_nm10_ & new_n_n15_;
  assign new_n_n45_ = new_nh10_ & new_ne10_ & new_nk10_ & new_nd2_;
  assign new_na10_ = new_nh10_ & new_n_n12_ & new_n_n9_;
  assign new_nf10_ = new_nh10_ & new_ni10_;
  assign new_n_n63_ = new_n_n13_ & new_nd10_ & new_nc2_ & new_nq0_ & new_ny1_;
  assign new_n_n52_ = new_nl10_ & new_n_n15_;
  assign new_nt4_ = new_nf10_ & new_nf2_;
  assign new_nz9_ = new_n_n39_ | new_n_n40_;
  assign new_ne10_ = new_n_n18_ & new_n_n22_ & new_nv10_;
  assign new_n_n64_ = new_nc2_ & new_nd10_ & new_n_n7_ & new_nc10_;
  assign new_n_n51_ = new_n_n15_ & new_n_n7_ & new_nk10_ & new_nd10_;
  assign new_n_n44_ = new_nf10_ & new_ne2_;
  assign new_n_n40_ = new_na10_ & new_nh2_ & new_nr10_ & new_n_n19_;
  assign new_n_n35_ = new_n_n22_ & new_ne2_;
  assign new_n_n0_ = ~new_np1_;
  assign new_n_n65_ = new_nc2_ & new_nd10_ & new_n_n21_ & new_nc10_;
  assign new_n_n30_ = new_nk10_ & new_n_n16_;
  assign new_nr10_ = new_n_n27_ | new_nv10_;
  assign new_n_n21_ = ~new_nd2_;
  assign new_n_n10_ = ~new_nb2_;
  assign new_n_n66_ = new_nc2_ & new_n_n16_ & new_nz1_ & new_nc10_;
  assign new_nj10_ = new_n_n10_ & new_na2_;
  assign new_nq10_ = new_n_n16_ & new_nc2_ & new_nj10_ & new_n_n15_;
  assign new_n_n20_ = ~new_ns0_;
  assign new_n_n11_ = ~new_nc2_;
  assign new_nk10_ = new_nb2_ & new_n_n13_;
  assign new_ns10_ = new_n_n25_ | new_n_n26_;
  assign new_n_n23_ = ~new_nf2_;
  assign new_n_n12_ = ~new_nf_;
  assign new_nl10_ = new_n_n11_ & new_nb2_;
  assign new_n_n27_ = new_nf2_ & new_ne2_;
  assign new_n_n22_ = ~new_nh2_;
  assign new_n_n13_ = ~new_na2_;
  assign new_nu4_ = new_n_n42_ | new_n_n43_;
  assign new_n_n38_ = new_ns10_ & new_n_n22_;
  assign new_nh10_ = new_nc2_ & new_n_n15_;
  assign new_nn10_ = new_nb2_ & new_nf_;
  assign new_nv10_ = new_n_n23_ & new_n_n24_;
  assign new_n_n14_ = ~new_nb1_;
  assign new_n_n43_ = new_nf10_ & new_ng2_;
  assign new_nb10_ = new_n_n37_ | new_n_n38_;
  assign new_ni10_ = new_n_n32_ | new_n_n31_ | new_n_n30_;
  assign new_n_n28_ = new_n_n11_ & new_n_n12_;
  assign new_n_n24_ = ~new_ne2_;
  assign new_n_n15_ = ~new_nb_;
  assign new_n_n58_ = new_n_n15_ & new_np0_ & new_n_n11_ & new_n_n19_ & new_nj10_;
  assign new_n_n49_ = new_n_n15_ & new_n_n7_ & new_nd10_ & new_nc2_ & new_nj10_;
  assign new_n_n32_ = new_n_n12_ & new_n_n9_;
  assign new_np10_ = new_n_n14_ & new_nl10_ & new_n_n15_ & new_nf_ & new_n_n13_;
  assign new_nt10_ = new_n_n19_ & new_na2_ & new_nu10_;
  assign new_n_n16_ = ~new_nd10_;
  assign new_n_n57_ = new_nn10_ & new_na2_ & new_nh10_ & new_n_n19_ & new_n_n6_;
  assign new_n_n50_ = new_n_n15_ & new_n_n21_ & new_nk10_ & new_nd10_;
  assign new_n_n31_ = new_nj10_ & new_n_n16_;
  assign new_no10_ = new_nl2_ & new_nf_ & new_n_n13_;
  assign new_nu10_ = new_n_n24_ | new_n_n23_ | new_nx1_ | new_n_n21_ | new_n_n22_ | new_n_n20_ | new_ng2_;
  assign new_n_n17_ = ~new_nr10_;
  assign new_n_n59_ = new_nn10_ & new_na2_ & new_nh10_ & new_n_n5_ & new_nr0_;
  assign new_np4_ = new_n_n54_ | new_n_n56_ | new_n_n55_ | new_n_n53_;
  assign new_nr4_ = new_n_n47_ | new_n_n46_ | new_n_n45_;
  assign new_ny9_ = new_n_n41_ | new_nz9_;
  assign new_n_n36_ = new_nh2_ & new_n_n24_;
  assign new_n_n26_ = new_nr10_ & new_ng2_;
  assign new_n_n18_ = ~new_ng2_;
  assign new_n_n60_ = new_n_n15_ & new_n_n11_ & new_nk10_;
  assign new_n_n56_ = new_n_n15_ & new_na2_ & new_nl10_;
  assign new_n_n48_ = new_n_n15_ & new_n_n21_ & new_nd10_ & new_nc2_ & new_nj10_;
  assign new_n_n41_ = new_na10_ & new_nb10_ & new_nr0_;
  assign new_nd10_ = new_n_n35_ | new_n_n36_;
  assign new_n_n25_ = new_n_n17_ & new_n_n18_;
  assign new_n_n19_ = ~new_nr0_;
  assign new_n_n61_ = new_n_n15_ & new_n_n11_ & new_n_n12_;
  assign new_n_n55_ = new_n_n15_ & new_np0_ & new_n_n11_ & new_na2_;
  assign new_n_n46_ = new_nh10_ & new_ne10_ & new_nj10_ & new_nd2_;
  assign new_n_n42_ = new_n_n15_ & new_nf_ & new_n_n13_ & new_nl10_;
  assign new_nc10_ = new_n_n10_ | new_n_n13_;
  assign new_n_n34_ = new_nn10_ & new_n_n15_ & new_n_n11_;
  assign new_n_n29_ = new_nn10_ & new_nt10_;
  assign new_no4_ = new_n_n59_ | new_n_n61_ | new_n_n60_ | new_n_n58_ | new_n_n57_;
  assign new_n_n54_ = new_n_n15_ & new_np0_ & new_nn10_ & new_na2_;
  assign new_n_n47_ = new_nh10_ & new_nd2_ & new_ni10_;
  assign new_nv4_ = new_nf10_ & new_nh2_;
  assign new_n_n37_ = new_n_n8_ & new_nh2_;
  assign new_n_n33_ = new_nn10_ & new_n_n15_ & new_nt10_;
  assign new_nm10_ = new_n_n28_ | new_n_n29_;
endmodule


