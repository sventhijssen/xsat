// Benchmark "parity" written by ABC on Sat Apr 29 10:30:09 2023

module parity ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
    f0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15;
  output f0;
  assign f0 = ((x14 ^ x15) & (((~x12 ^ x13) & (((~x10 ^ x11) & (((~x8 ^ x9) & (((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))) | ((x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))))) | ((x10 ^ x11) & (((((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))) & (x8 ^ x9)) | ((~x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))))))) | ((x12 ^ x13) & (((((~x8 ^ x9) & (((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))) | ((x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))))) & (x10 ^ x11)) | ((~x10 ^ x11) & (((((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))) & (x8 ^ x9)) | ((~x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))))))))) | ((~x14 ^ x15) & (((((~x10 ^ x11) & (((~x8 ^ x9) & (((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))) | ((x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))))) | ((x10 ^ x11) & (((((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))) & (x8 ^ x9)) | ((~x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))))))) & (x12 ^ x13)) | ((~x12 ^ x13) & (((((~x8 ^ x9) & (((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))))) | ((x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))))) & (x10 ^ x11)) | ((~x10 ^ x11) & (((((~x6 ^ x7) & (((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1)))))) | ((x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))) & (x8 ^ x9)) | ((~x8 ^ x9) & (((((~x4 ^ x5) & (((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1)))) | ((x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))) & (x6 ^ x7)) | ((~x6 ^ x7) & (((((~x2 ^ x3) & (~x0 ^ x1)) | ((x2 ^ x3) & (x0 ^ x1))) & (x4 ^ x5)) | ((~x4 ^ x5) & (((~x0 ^ x1) & (x2 ^ x3)) | ((~x2 ^ x3) & (x0 ^ x1))))))))))))));
endmodule


