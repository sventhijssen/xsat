// Benchmark "top" written by ABC on Fri Mar 31 12:11:47 2023

module top ( 
    pina0, pinb1, pinc2, pind3, pina1, pinb0, pinc3, pind2, pmusel1, pinc4,
    pind5, pmusel2, pinc5, pind4, pmusel3, pina4, pinb5, pina5, pinb4,
    pina2, pinb3, pinc0, pind1, pina3, pinb2, pinc1, pind0, pind15, pinc15,
    pind14, pinb15, pinc14, pind13, popsel3, popsel1, popsel2, pina11,
    pinb10, pina10, popsel0, pina15, pinb14, pinc13, pind12, pina14,
    pinb13, pinc12, pind11, pina13, pinb12, pinc11, pind10, pina12, pinb11,
    pinc10, pina8, pinb9, pina9, pinb8, pina6, pinb7, pina7, pinb6, psh0,
    pinc6, pind7, pmusel4, psh1, pinc7, pind6, psh2, pinc8, pind9, pinc9,
    pind8,
    po12, po11, po14, po13, po15, po9, po8, po7, po6, po5, po4, po3, po2,
    po1, po0, po10  );
  input  pina0, pinb1, pinc2, pind3, pina1, pinb0, pinc3, pind2, pmusel1,
    pinc4, pind5, pmusel2, pinc5, pind4, pmusel3, pina4, pinb5, pina5,
    pinb4, pina2, pinb3, pinc0, pind1, pina3, pinb2, pinc1, pind0, pind15,
    pinc15, pind14, pinb15, pinc14, pind13, popsel3, popsel1, popsel2,
    pina11, pinb10, pina10, popsel0, pina15, pinb14, pinc13, pind12,
    pina14, pinb13, pinc12, pind11, pina13, pinb12, pinc11, pind10, pina12,
    pinb11, pinc10, pina8, pinb9, pina9, pinb8, pina6, pinb7, pina7, pinb6,
    psh0, pinc6, pind7, pmusel4, psh1, pinc7, pind6, psh2, pinc8, pind9,
    pinc9, pind8;
  output po12, po11, po14, po13, po15, po9, po8, po7, po6, po5, po4, po3, po2,
    po1, po0, po10;
  wire new_nina0_, new_ninb1_, new_ninc2_, new_nind3_, new_nina1_,
    new_ninb0_, new_ninc3_, new_nind2_, new_nmusel1_, new_ninc4_,
    new_nind5_, new_nmusel2_, new_ninc5_, new_nind4_, new_nmusel3_,
    new_nina4_, new_ninb5_, new_nina5_, new_ninb4_, new_nina2_, new_ninb3_,
    new_ninc0_, new_nind1_, new_nina3_, new_ninb2_, new_ninc1_, new_nind0_,
    new_nind15_, new_ninc15_, new_nind14_, new_ninb15_, new_ninc14_,
    new_nind13_, new_nopsel3_, new_nopsel1_, new_nopsel2_, new_nina11_,
    new_ninb10_, new_nina10_, new_nopsel0_, new_nina15_, new_ninb14_,
    new_ninc13_, new_nind12_, new_nina14_, new_ninb13_, new_ninc12_,
    new_nind11_, new_nina13_, new_ninb12_, new_ninc11_, new_nind10_,
    new_nina12_, new_ninb11_, new_ninc10_, new_nina8_, new_ninb9_,
    new_nina9_, new_ninb8_, new_nina6_, new_ninb7_, new_nina7_, new_ninb6_,
    new_nsh0_, new_ninc6_, new_nind7_, new_nmusel4_, new_nsh1_, new_ninc7_,
    new_nind6_, new_nsh2_, new_ninc8_, new_nind9_, new_ninc9_, new_nind8_,
    new_n_n2456_, new_n_n1583_, new_n_n2439_, new_n_n2385_, new_n_n2380_,
    new_n_n2372_, new_n_n1546_, new_n_n1542_, new_n_n1536_, new_n_n1517_,
    new_n_n2329_, new_n_n1508_, new_n_n2317_, new_n_n2312_, new_n_n1493_,
    new_n_n1486_, new_n_n2297_, new_n_n2291_, new_n_n1460_, new_n_n2271_,
    new_n_n2265_, new_n_n1446_, new_n_n2255_, new_n_n2247_, new_n_n1430_,
    new_n_n1424_, new_n_n1398_, new_n_n2208_, new_n_n2200_, new_n_n1383_,
    new_n_n2190_, new_n_n1330_, new_n_n1956_, new_n_n1953_, new_n_n1064_,
    new_n_n1907_, new_n_n1900_, new_n_n1896_, new_n_n1891_, new_n_n1868_,
    new_n_n1011_, new_n_n1858_, new_n_n1855_, new_n_n990_, new_n_n985_,
    new_n_n1841_, new_n_n1836_, new_n_n960_, new_n_n955_, new_n_n1809_,
    new_n_n943_, new_n_n937_, new_n_n1795_, new_n_n1790_, new_n_n1785_,
    new_n_n914_, new_n_n890_, new_n_n886_, new_n_n879_, new_n_n871_,
    new_ne0_, new_n_n1740_, new_n_n858_, new_n_n851_, new_n_n1725_,
    new_n_n838_, new_n_n1718_, new_n_n1716_, new_n_n785_, new_n_n775_,
    new_n_n767_, new_n_n758_, new_n_n748_, new_n_n737_, new_n_n1699_,
    new_n_n1692_, new_n_n696_, new_n_n686_, new_n_n676_, new_n_n668_,
    new_n_n1680_, new_n_n648_, new_n_n640_, new_n_n622_, new_n_n611_,
    new_n_n601_, new_n_n594_, new_n_n585_, new_n_n575_, new_n_n567_,
    new_n_n1660_, new_n_n548_, new_n_n540_, new_n_n531_, new_n_n521_,
    new_n_n510_, new_n_n501_, new_n_n492_, new_n_n482_, new_n_n471_,
    new_n_n462_, new_n_n452_, new_n_n442_, new_n_n434_, new_n_n427_,
    new_n_n419_, new_n_n1633_, new_n_n400_, new_n_n391_, new_n_n380_,
    new_n_n372_, new_n_n354_, new_n_n344_, new_n_n1620_, new_n_n327_,
    new_n_n317_, new_n_n1614_, new_n_n296_, new_n_n286_, new_n_n256_,
    new_n_n245_, new_n_n235_, new_n_n225_, new_n_n215_, new_n_n204_,
    new_n_n194_, new_n_n153_, new_n_n1602_, new_n_n132_, new_n_n122_,
    new_n_n112_, new_n_n101_, new_n_n1586_, new_n_n2447_, new_n_n2440_,
    new_n_n1561_, new_n_n2379_, new_n_n2373_, new_n_n2367_, new_n_n2362_,
    new_n_n1532_, new_n_n1518_, new_n_n2328_, new_n_n2323_, new_nb3_,
    new_n_n2313_, new_n_n1492_, new_n_n1487_, new_n_n1480_, new_nb1_,
    new_n_n1466_, new_n_n2270_, new_n_n2266_, new_n_n1445_, new_n_n1440_,
    new_n_n1436_, new_n_n1431_, new_n_n1423_, new_n_n2213_, new_n_n1393_,
    new_n_n1389_, new_n_n1384_, new_n_n2189_, new_ng3_, new_n_n1115_,
    new_n_n1109_, new_n_n1913_, new_n_n1908_, new_n_n1899_, new_n_n1050_,
    new_n_n1886_, new_n_n1867_, new_n_n1012_, new_n_n1004_, new_n_n997_,
    new_n_n1851_, new_n_n1846_, new_n_n978_, new_n_n973_, new_n_n965_,
    new_n_n954_, new_n_n1810_, new_n_n1803_, new_n_n1799_, new_no2_,
    new_n_n926_, new_n_n919_, new_n_n1780_, new_n_n1763_, new_n_n887_,
    new_n_n878_, new_n_n872_, new_n_n865_, new_n_n1741_, new_n_n1733_,
    new_n_n852_, new_n_n844_, new_n_n1721_, new_n_n829_, new_n_n1717_,
    new_n_n784_, new_n_n776_, new_n_n766_, new_n_n1702_, new_n_n747_,
    new_n_n738_, new_n_n721_, new_n_n701_, new_n_n1687_, new_n_n1685_,
    new_n_n677_, new_n_n667_, new_n_n659_, new_n_n647_, new_n_n641_,
    new_n_n621_, new_n_n612_, new_n_n600_, new_n_n595_, new_n_n584_,
    new_n_n576_, new_n_n566_, new_n_n558_, new_n_n541_, new_n_n539_,
    new_n_n532_, new_n_n520_, new_n_n511_, new_n_n500_, new_n_n1649_,
    new_n_n481_, new_n_n472_, new_n_n461_, new_n_n453_, new_n_n451_,
    new_n_n433_, new_n_n428_, new_n_n418_, new_n_n409_, new_n_n399_,
    new_n_n392_, new_n_n379_, new_n_n373_, new_n_n353_, new_n_n345_,
    new_n_n1619_, new_n_n1616_, new_n_n316_, new_n_n307_, new_n_n295_,
    new_n_n287_, new_n_n265_, new_n_n244_, new_n_n236_, new_n_n224_,
    new_n_n216_, new_n_n203_, new_n_n1606_, new_n_n152_, new_n_n143_,
    new_n_n131_, new_n_n123_, new_n_n111_, new_n_n102_, new_n_n2454_,
    new_n_n2449_, new_n_n2441_, new_n_n1560_, new_n_n1556_, new_n_n2374_,
    new_n_n2366_, new_n_n2357_, new_n_n1533_, new_n_n2335_, new_n_n1513_,
    new_n_n2324_, new_n_n2316_, new_n_n1497_, new_n_n2306_, new_n_n1488_,
    new_n_n2287_, new_n_n1471_, new_n_n1455_, new_n_n1450_, new_n_n2259_,
    new_n_n1441_, new_n_n1435_, new_n_n1428_, new_n_n2240_, new_n_n1409_,
    new_n_n1402_, new_n_n1388_, new_n_n2196_, new_n_n1379_, new_n_n2155_,
    new_n_n1169_, new_n_n1958_, new_n_n1110_, new_n_n1914_, new_n_n1909_,
    new_n_n1898_, new_n_n1892_, new_n_n1887_, new_n_n1018_, new_n_n1013_,
    new_n_n1003_, new_n_n995_, new_no4_, new_n_n1847_, new_n_n1831_,
    new_n_n966_, new_n_n953_, new_n_n948_, new_n_n1804_, new_n_n938_,
    new_n_n930_, new_n_n925_, new_n_n920_, new_n_n915_, new_n_n1770_,
    new_n_n1767_, new_n_n877_, new_n_n1749_, new_n_n866_, new_n_n1742_,
    new_n_n859_, new_n_n853_, new_n_n843_, new_n_n836_, new_n_n1719_,
    new_n_n821_, new_n_n787_, new_n_n777_, new_n_n1703_, new_n_n756_,
    new_n_n750_, new_n_n739_, new_n_n712_, new_n_n1693_, new_n_n1688_,
    new_n_n685_, new_n_n1684_, new_n_n670_, new_n_n660_, new_n_n633_,
    new_n_n623_, new_n_n613_, new_n_n1671_, new_n_n593_, new_n_n1666_,
    new_n_n577_, new_n_n565_, new_n_n550_, new_n_n542_, new_n_n519_,
    new_n_n508_, new_n_n502_, new_n_n493_, new_n_n480_, new_n_n469_,
    new_n_n464_, new_n_n454_, new_n_n432_, new_n_n425_, new_n_n420_,
    new_n_n410_, new_n_n398_, new_n_n389_, new_n_n382_, new_n_n1626_,
    new_n_n352_, new_n_n342_, new_n_n335_, new_n_n328_, new_n_n315_,
    new_n_n305_, new_n_n298_, new_n_n288_, new_n_n264_, new_n_n254_,
    new_n_n237_, new_n_n223_, new_n_n213_, new_n_n206_, new_n_n195_,
    new_n_n171_, new_n_n161_, new_n_n130_, new_n_n120_, new_n_n114_,
    new_n_n103_, new_n_n2455_, new_n_n2448_, new_n_n1581_, new_n_n2384_,
    new_n_n1555_, new_n_n2375_, new_n_n1541_, new_n_n1537_, new_n_n1534_,
    new_n_n1516_, new_n_n2330_, new_n_n2325_, new_n_n1502_, new_n_n2311_,
    new_n_n1494_, new_n_n1489_, new_n_n2286_, new_n_n2269_, new_n_n2264_,
    new_n_n1447_, new_n_n1442_, new_n_n1434_, new_n_n1429_, new_n_n2239_,
    new_n_n1408_, new_n_n1403_, new_n_n1387_, new_n_n1382_, new_n_n2191_,
    new_n_n2159_, new_n_n1994_, new_n_n1957_, new_n_n1111_, new_n_n1065_,
    new_n_n1060_, new_no6_, new_n_n1045_, new_n_n1040_, new_n_n1017_,
    new_n_n1863_, new_n_n1857_, new_n_n996_, new_n_n991_, new_n_n986_,
    new_n_n1830_, new_ne3_, new_n_n1813_, new_n_n1808_, new_n_n944_,
    new_n_n939_, new_n_n1794_, new_n_n1789_, new_n_n1786_, new_n_n1781_,
    new_n_n902_, new_n_n896_, new_n_n1752_, new_n_n870_, new_n_n1745_,
    new_n_n861_, new_n_n1734_, new_n_n854_, new_n_n842_, new_n_n837_,
    new_n_n830_, new_n_n822_, new_n_n786_, new_n_n778_, new_n_n765_,
    new_n_n757_, new_n_n749_, new_n_n740_, new_n_n703_, new_n_n702_,
    new_n_n1689_, new_n_n684_, new_n_n675_, new_n_n669_, new_n_n661_,
    new_n_n632_, new_n_n624_, new_n_n1673_, new_n_n599_, new_n_n1667_,
    new_n_n586_, new_n_n578_, new_n_n557_, new_n_n549_, new_n_n1656_,
    new_n_n518_, new_n_n509_, new_n_n1651_, new_n_n494_, new_n_n479_,
    new_n_n470_, new_n_n463_, new_n_n455_, new_n_n1640_, new_n_n426_,
    new_n_n1634_, new_n_n411_, new_n_n397_, new_n_n390_, new_n_n381_,
    new_n_n1627_, new_n_n351_, new_n_n343_, new_n_n334_, new_n_n329_,
    new_n_n314_, new_n_n306_, new_n_n297_, new_n_n289_, new_n_n263_,
    new_n_n255_, new_n_n246_, new_n_n222_, new_n_n214_, new_n_n205_,
    new_n_n196_, new_n_n170_, new_n_n162_, new_n_n1601_, new_n_n121_,
    new_n_n113_, new_n_n104_, new_n_n2459_, new_n_n1584_, new_n_n2442_,
    new_n_n1562_, new_n_n2381_, new_n_n1552_, new_n_n1528_, new_n_n2341_,
    new_n_n2336_, new_n_n1501_, new_n_n2310_, new_n_n2299_, new_n_n1478_,
    new_n_n2289_, new_n_n1454_, new_n_n2263_, new_n_n2257_, new_n_n1439_,
    new_n_n1437_, new_n_n1433_, new_n_n2242_, new_n_n2221_, new_n_n2217_,
    new_n_n1397_, new_n_n1392_, new_n_n1380_, new_n_n2163_, new_n_n2000_,
    new_n_n1165_, new_n_n1117_, new_n_n1954_, new_n_n1067_, new_n_n1061_,
    new_n_n1882_, new_n_n1877_, new_n_n1024_, new_n_n1002_, new_n_n1854_,
    new_n_n1843_, new_n_n1837_, new_n_n969_, new_n_n967_, new_n_n1812_,
    new_n_n947_, new_n_n941_, new_n_n935_, new_n_n933_, new_n_n927_,
    new_n_n922_, new_n_n1782_, new_n_n901_, new_n_n1765_, new_n_n1760_,
    new_n_n883_, new_n_n1746_, new_no0_, new_n_n1731_, new_n_n849_,
    new_n_n846_, new_n_n1722_, new_n_n832_, new_n_n823_, new_n_n782_,
    new_n_n771_, new_n_n1705_, new_n_n761_, new_n_n752_, new_n_n741_,
    new_n_n699_, new_n_n692_, new_n_n690_, new_n_n680_, new_n_n671_,
    new_n_n662_, new_n_n618_, new_n_n608_, new_n_n1668_, new_n_n588_,
    new_n_n579_, new_n_n537_, new_n_n528_, new_n_n504_, new_n_n1650_,
    new_n_n448_, new_n_n438_, new_n_n412_, new_n_n396_, new_n_n369_,
    new_n_n360_, new_n_n313_, new_n_n303_, new_n_n282_, new_n_n273_,
    new_n_n221_, new_n_n211_, new_n_n200_, new_n_n190_, new_n_n180_,
    new_n_n129_, new_n_n118_, new_n_n108_, new_n_n97_, new_n_n8_,
    new_n_n1587_, new_n_n2450_, new_n_n2443_, new_n_n1557_, new_n_n2376_,
    new_n_n1527_, new_n_n2342_, new_n_n2315_, new_n_n1496_, new_n_n2298_,
    new_n_n1479_, new_n_n2288_, new_n_n2268_, new_n_n1449_, new_n_n1444_,
    new_n_n2252_, new_n_n2250_, new_n_n2245_, new_n_n2241_, new_nb4_,
    new_n_n2218_, new_n_n2210_, new_n_n2205_, new_n_n2192_, new_n_n2170_,
    new_n_n1170_, new_n_n1995_, new_n_n1116_, new_n_n1955_, new_n_n1066_,
    new_n_n1062_, new_n_n1035_, new_n_n1030_, new_n_n1019_, new_n_n1001_,
    new_n_n994_, new_n_n1842_, new_n_n976_, new_n_n1832_, new_n_n968_,
    new_n_n952_, new_n_n1807_, new_n_n1801_, new_n_n936_, new_n_n1796_,
    new_n_n928_, new_n_n921_, new_n_n1783_, new_n_n900_, new_n_n1766_,
    new_n_n889_, new_n_n884_, new_n_n867_, new_n_n1743_, new_n_n856_,
    new_n_n1728_, new_n_n1727_, new_n_n1723_, new_n_n831_, new_n_n824_,
    new_n_n781_, new_n_n772_, new_n_n1704_, new_n_n762_, new_n_n751_,
    new_n_n742_, new_n_n698_, new_n_n693_, new_n_n689_, new_n_n681_,
    new_n_n1682_, new_n_n663_, new_n_n617_, new_n_n609_, new_n_n604_,
    new_n_n587_, new_n_n580_, new_n_n536_, new_n_n1653_, new_n_n503_,
    new_n_n495_, new_n_n447_, new_n_n439_, new_n_n421_, new_n_n388_,
    new_n_n368_, new_n_n1623_, new_n_n312_, new_n_n304_, new_n_n281_,
    new_n_n1611_, new_n_n220_, new_n_n212_, new_n_n191_, new_n_n189_,
    new_n_n181_, new_n_n128_, new_n_n119_, new_n_n107_, new_n_n98_,
    new_n_n2457_, new_n_n2452_, new_n_n2444_, new_n_n2386_, new_n_n1553_,
    new_n_n2347_, new_n_n1520_, new_n_n2305_, new_n_n1485_, new_n_n1482_,
    new_n_n2292_, new_n_n1473_, new_n_n1453_, new_n_n2262_, new_n_n2258_,
    new_n_n2253_, new_n_n2249_, new_n_n2244_, new_n_n1426_, new_n_n2220_,
    new_n_n2215_, new_n_n2212_, new_n_n2206_, new_n_n2202_, new_n_n2197_,
    new_nb9_, new_n_n2050_, new_n_n2043_, new_n_n1171_, new_n_n1166_,
    new_n_n1959_, new_n_n1112_, new_n_n1910_, new_n_n1881_, new_n_n1025_,
    new_n_n1869_, new_n_n1850_, new_n_n984_, new_n_n980_, new_n_n974_,
    new_n_n1833_, new_n_n1824_, new_n_n951_, new_n_n945_, new_n_n1802_,
    new_n_n1797_, new_n_n932_, new_n_n1791_, new_n_n923_, new_n_n916_,
    new_n_n899_, new_n_n894_, new_n_n1762_, new_n_n885_, new_n_n1753_,
    new_n_n1750_, new_n_n857_, new_n_n1729_, new_n_n1726_, new_n_n839_,
    new_n_n834_, new_n_n825_, new_n_n783_, new_n_n773_, new_n_n769_,
    new_n_n759_, new_n_n753_, new_n_n743_, new_n_n700_, new_n_n694_,
    new_n_n688_, new_n_n678_, new_n_n673_, new_n_n1681_, new_n_n620_,
    new_n_n610_, new_n_n603_, new_n_n596_, new_n_n581_, new_n_n1655_,
    new_n_n529_, new_n_n523_, new_n_n512_, new_n_n450_, new_n_n440_,
    new_n_n429_, new_n_n378_, new_n_n1625_, new_n_n361_, new_n_n294_,
    new_n_n284_, new_n_n274_, new_n_n219_, new_n_n202_, new_n_n192_,
    new_n_n127_, new_n_n1600_, new_n_n110_, new_n_n99_, new_n_n2458_,
    new_n_n2451_, new_n_n1582_, new_n_n2387_, new_n_n1558_, new_n_n2340_,
    new_n_n1519_, new_nb2_, new_n_n2302_, new_n_n1481_, new_n_n1477_,
    new_n_n1472_, new_n_n1452_, new_n_n1448_, new_nb7_, new_n_n2254_,
    new_n_n2248_, new_n_n1432_, new_n_n1425_, new_n_n1407_, new_n_n2216_,
    new_n_n2211_, new_n_n2207_, new_n_n2201_, new_n_n1385_, new_n_n2179_,
    new_n_n2049_, new_n_n2044_, new_n_n2001_, new_n_n1996_, new_n_n1118_,
    new_n_n1113_, new_n_n1915_, new_n_n1876_, new_ne5_, new_n_n1870_,
    new_n_n989_, new_n_n1845_, new_n_n979_, new_n_n975_, new_n_n970_,
    new_n_n1825_, new_n_n1811_, new_n_n946_, new_n_n942_, new_n_n1798_,
    new_n_n931_, new_n_n1792_, new_n_n1787_, new_n_n917_, new_n_n1769_,
    new_n_n895_, new_n_n1761_, new_n_n1756_, new_n_n880_, new_n_n873_,
    new_n_n1732_, new_n_n850_, new_n_n845_, new_n_n840_, new_n_n833_,
    new_n_n826_, new_n_n1707_, new_n_n774_, new_n_n768_, new_n_n760_,
    new_n_n1701_, new_n_n744_, new_n_n1691_, new_n_n695_, new_n_n687_,
    new_n_n679_, new_n_n672_, new_n_n664_, new_n_n619_, new_n_n1672_,
    new_n_n602_, new_n_n597_, new_n_n589_, new_n_n538_, new_n_n530_,
    new_n_n522_, new_n_n513_, new_n_n449_, new_n_n441_, new_n_n1641_,
    new_n_n371_, new_n_n370_, new_n_n362_, new_n_n1613_, new_n_n285_,
    new_n_n283_, new_n_n210_, new_n_n201_, new_n_n193_, new_n_n126_,
    new_n_n117_, new_n_n109_, new_n_n100_, new_n_n2484_, new_n_n2477_,
    new_n_n2437_, new_n_n1577_, new_n_n2420_, new_n_n2412_, new_n_n1569_,
    new_n_n2395_, new_n_n1564_, new_n_n2365_, new_n_n1540_, new_n_n2355_,
    new_n_n1531_, new_n_n1525_, new_nb12_, new_n_n2331_, new_n_n1484_,
    new_n_n2295_, new_n_n2290_, new_n_n2282_, new_n_n1463_, new_n_n1457_,
    new_n_n2235_, new_n_n1416_, new_n_n2225_, new_n_n2184_, new_n_n2038_,
    new_n_n1201_, new_n_n1992_, new_n_n1155_, new_n_n1982_, new_n_n1978_,
    new_n_n1973_, new_n_n1951_, new_n_n1102_, new_n_n1096_, new_n_n1935_,
    new_n_n1085_, new_n_n1079_, new_n_n1921_, new_n_n1916_, new_n_n1055_,
    new_n_n1895_, new_n_n1889_, new_n_n1037_, new_n_n1879_, new_n_n1873_,
    new_n_n1020_, new_n_n1844_, new_n_n1840_, new_n_n972_, new_n_n1826_,
    new_n_n1821_, new_n_n1815_, new_n_n1784_, new_n_n1777_, new_n_n906_,
    new_n_n1714_, new_n_n810_, new_n_n1711_, new_n_n792_, new_n_n735_,
    new_n_n727_, new_n_n717_, new_n_n708_, new_n_n656_, new_n_n645_,
    new_n_n638_, new_n_n628_, new_n_n614_, new_n_n1661_, new_n_n555_,
    new_n_n545_, new_n_n533_, new_n_n524_, new_n_n468_, new_n_n460_,
    new_n_n445_, new_n_n436_, new_n_n430_, new_n_n377_, new_n_n366_,
    new_n_n357_, new_n_n1621_, new_n_n336_, new_n_n279_, new_n_n269_,
    new_n_n258_, new_n_n248_, new_n_n238_, new_n_n186_, new_n_n176_,
    new_n_n166_, new_n_n1603_, new_n_n145_, new_n_n135_, new_n_n5_,
    new_n_n2485_, new_n_n2469_, new_n_n2436_, new_n_n2429_, new_n_n1574_,
    new_n_n1572_, new_n_n2403_, new_n_n2396_, new_n_n1563_, new_n_n2371_,
    new_n_n1539_, new_n_n1535_, new_n_n1530_, new_n_n1526_, new_n_n2337_,
    new_n_n1514_, new_n_n1483_, new_n_n2296_, new_n_n1474_, new_n_n2283_,
    new_n_n1462_, new_n_n2273_, new_n_n1427_, new_n_n2236_, new_n_n1415_,
    new_n_n1411_, new_n_n2187_, new_n_n1207_, new_n_n1202_, new_n_n1160_,
    new_n_n1987_, new_n_n1981_, new_n_n1143_, new_n_n1968_, new_n_n1950_,
    new_n_n1946_, new_n_n1095_, new_n_n1936_, new_n_n1929_, new_n_n1926_,
    new_n_n1073_, new_n_n1068_, new_n_n1905_, new_n_n1894_, new_n_n1044_,
    new_n_n1036_, new_n_n1880_, new_n_n1026_, new_no5_, new_n_n983_,
    new_n_n977_, new_n_n971_, new_n_n1827_, new_n_n1820_, new_n_n957_,
    new_n_n924_, new_n_n910_, new_n_n1771_, new_n_n1713_, new_n_n811_,
    new_n_n800_, new_n_n793_, new_n_n734_, new_n_n1697_, new_n_n1695_,
    new_n_n709_, new_n_n655_, new_n_n646_, new_n_n637_, new_n_n629_,
    new_n_n605_, new_n_n1664_, new_n_n554_, new_n_n546_, new_n_n1654_,
    new_n_n525_, new_n_n1647_, new_n_n1645_, new_n_n444_, new_n_n1642_,
    new_n_n1635_, new_n_n387_, new_n_n365_, new_n_n358_, new_n_n346_,
    new_n_n337_, new_n_n278_, new_n_n270_, new_n_n257_, new_n_n249_,
    new_n_n229_, new_n_n185_, new_n_n177_, new_n_n165_, new_n_n156_,
    new_n_n144_, new_n_n136_, new_n_n6_, new_n_n2486_, new_n_n2462_,
    new_n_n2435_, new_n_n2427_, new_n_n2422_, new_n_n2413_, new_n_n2402_,
    new_n_n2394_, new_n_n2389_, new_nb15_, new_n_n1545_, new_n_n2356_,
    new_n_n2348_, new_n_n1524_, new_n_n1521_, new_n_n1509_, new_n_n2319_,
    new_n_n2301_, new_n_n2293_, new_n_n1476_, new_n_n1468_, new_n_n1464_,
    new_n_n1458_, new_nb6_, new_n_n1421_, new_n_n1417_, new_n_n2226_,
    new_n_n1197_, new_n_n1191_, new_n_n1159_, new_n_n1153_, new_n_n1150_,
    new_n_n1144_, new_n_n1127_, new_n_n1107_, new_n_n1945_, new_n_n1941_,
    new_n_n1091_, new_n_n1084_, new_n_n1925_, new_n_n1074_, new_n_n1069_,
    new_n_n1904_, new_ne6_, new_n_n1890_, new_n_n1884_, new_n_n1031_,
    new_n_n1027_, new_n_n1871_, new_n_n1864_, new_n_n1008_, new_n_n982_,
    new_n_n1838_, new_n_n1835_, new_n_n1828_, new_no3_, new_n_n1816_,
    new_n_n929_, new_n_n1779_, new_n_n1772_, new_n_n819_, new_n_n808_,
    new_n_n801_, new_n_n794_, new_n_n780_, new_n_n733_, new_n_n725_,
    new_n_n719_, new_n_n710_, new_n_n1690_, new_n_n1686_, new_n_n654_,
    new_n_n644_, new_n_n639_, new_n_n630_, new_n_n616_, new_n_n606_,
    new_n_n571_, new_n_n563_, new_n_n547_, new_n_n535_, new_n_n526_,
    new_n_n488_, new_n_n477_, new_n_n1644_, new_n_n437_, new_n_n413_,
    new_n_n1630_, new_n_n367_, new_n_n1622_, new_n_n330_, new_n_n321_,
    new_n_n1612_, new_n_n271_, new_n_n1610_, new_n_n240_, new_n_n230_,
    new_n_n188_, new_n_n178_, new_n_n164_, new_n_n154_, new_n_n147_,
    new_n_n137_, new_n_n1597_, new_n_n1579_, new_n_n2428_, new_n_n2421_,
    new_n_n2414_, new_n_n2401_, new_n_n1566_, new_n_n2388_, new_n_n2370_,
    new_n_n2364_, new_n_n2361_, new_n_n1529_, new_n_n2343_, new_n_n2338_,
    new_n_n2326_, new_n_n2320_, new_n_n2300_, new_n_n2294_, new_n_n1475_,
    new_n_n2281_, new_n_n2278_, new_n_n1459_, new_n_n2251_, new_n_n2234_,
    new_n_n2231_, new_n_n1412_, new_n_n1196_, new_n_n1192_, new_n_n1991_,
    new_n_n1154_, new_n_n1149_, new_n_n1979_, new_n_n1960_, new_n_n1949_,
    new_n_n1101_, new_n_n1097_, new_n_n1092_, new_n_n1928_, new_n_n1078_,
    new_n_n1922_, new_n_n1070_, new_n_n1903_, new_n_n1054_, new_n_n1049_,
    new_n_n1883_, new_n_n1878_, new_n_n1874_, new_n_n1021_, new_n_n1014_,
    new_n_n1860_, new_n_n981_, new_n_n1839_, new_n_n1834_, new_n_n1829_,
    new_n_n962_, new_n_n1817_, new_n_n934_, new_n_n1778_, new_n_n907_,
    new_n_n818_, new_n_n809_, new_n_n1712_, new_n_n795_, new_n_n770_,
    new_n_n732_, new_n_n726_, new_n_n718_, new_n_n711_, new_n_n697_,
    new_n_n691_, new_n_n653_, new_n_n1679_, new_n_n1676_, new_n_n631_,
    new_n_n615_, new_n_n607_, new_n_n1663_, new_n_n564_, new_n_n556_,
    new_n_n534_, new_n_n527_, new_n_n487_, new_n_n478_, new_n_n446_,
    new_n_n1643_, new_n_n405_, new_n_n1631_, new_n_n1624_, new_n_n359_,
    new_n_n1617_, new_n_n322_, new_n_n280_, new_n_n272_, new_n_n247_,
    new_n_n239_, new_n_n1608_, new_n_n187_, new_n_n179_, new_n_n163_,
    new_n_n155_, new_n_n146_, new_n_n138_, new_n_n7_, new_n_n2479_,
    new_n_n1591_, new_n_n2463_, new_n_n2434_, new_n_n1576_, new_n_n2417_,
    new_n_n2409_, new_n_n1570_, new_n_n2398_, new_npgx3_, new_n_n2382_,
    new_n_n1554_, new_n_n1548_, new_n_n1543_, new_n_n2359_, new_n_n2351_,
    new_n_n2346_, new_n_n1523_, new_n_n2333_, new_n_n1511_, new_n_n2321_,
    new_n_n2318_, new_n_n1499_, new_n_n2308_, new_n_n2303_, new_n_n2285_,
    new_n_n2279_, new_n_n2274_, new_n_n2256_, new_n_n2232_, new_n_n1413_,
    new_n_n2022_, new_n_n1181_, new_n_n1158_, new_n_n1139_, new_n_n1134_,
    new_n_n1128_, new_n_n1961_, new_n_n1106_, new_n_n1099_, new_n_n1938_,
    new_n_n1089_, new_n_n1931_, new_ne7_, new_n_n1076_, new_n_n1917_,
    new_n_n1063_, new_n_n1902_, new_n_n1052_, new_n_n1046_, new_n_n1041_,
    new_n_n1034_, new_n_n1875_, new_n_n1022_, new_n_n1865_, new_n_n1009_,
    new_n_n1007_, new_n_n999_, new_n_n993_, new_n_n1848_, new_n_n963_,
    new_n_n958_, new_n_n1800_, new_n_n912_, new_n_n908_, new_n_n817_,
    new_n_n806_, new_n_n798_, new_n_n1708_, new_n_n764_, new_n_n731_,
    new_n_n1696_, new_n_n714_, new_n_n704_, new_n_n683_, new_n_n674_,
    new_n_n652_, new_n_n642_, new_n_n1675_, new_n_n625_, new_n_n598_,
    new_n_n591_, new_n_n1665_, new_n_n1662_, new_n_n561_, new_n_n552_,
    new_n_n1657_, new_n_n517_, new_n_n506_, new_n_n497_, new_n_n489_,
    new_n_n486_, new_n_n475_, new_n_n465_, new_n_n456_, new_n_n431_,
    new_n_n423_, new_n_n415_, new_n_n406_, new_n_n404_, new_n_n394_,
    new_n_n384_, new_n_n374_, new_n_n350_, new_n_n340_, new_n_n331_,
    new_n_n323_, new_n_n320_, new_n_n310_, new_n_n300_, new_n_n290_,
    new_n_n275_, new_n_n262_, new_n_n252_, new_n_n242_, new_n_n231_,
    new_n_n218_, new_n_n208_, new_n_n197_, new_n_n182_, new_n_n172_,
    new_n_n169_, new_n_n159_, new_n_n149_, new_n_n139_, new_n_n116_,
    new_n_n105_, new_n_n1_, new_n_n2478_, new_n_n2472_, new_n_n1588_,
    new_n_n2433_, new_n_n2426_, new_n_n1573_, new_n_n1571_, new_n_n2406_,
    new_n_n2399_, new_n_n2390_, new_n_n2383_, new_n_n1549_, new_n_n1547_,
    new_n_n1544_, new_n_n2358_, new_n_n2352_, new_n_n2350_, new_n_n1522_,
    new_n_n2334_, new_n_n1510_, new_n_n1506_, new_n_n1505_, new_n_n1500_,
    new_n_n2307_, new_n_n1490_, new_n_n1470_, new_n_n1465_, new_n_n2275_,
    new_n_n2260_, new_n_n1418_, new_n_n2227_, new_n_n2021_, new_n_n2016_,
    new_n_n1986_, new_n_n1975_, new_n_n1135_, new_n_n1964_, new_n_n1121_,
    new_n_n1948_, new_n_n1100_, new_n_n1094_, new_n_n1933_, new_n_n1087_,
    new_n_n1082_, new_n_n1075_, new_n_n1071_, new_n_n1906_, new_n_n1901_,
    new_n_n1053_, new_n_n1893_, new_n_n1042_, new_n_n1039_, new_n_n1028_,
    new_n_n1872_, new_n_n1015_, new_n_n1010_, new_n_n1859_, new_n_n1000_,
    new_n_n992_, new_n_n1849_, new_n_n1822_, new_n_n1818_, new_n_n1805_,
    new_n_n911_, new_n_n1773_, new_n_n816_, new_n_n807_, new_n_n797_,
    new_n_n789_, new_n_n755_, new_n_n730_, new_n_n724_, new_n_n713_,
    new_n_n705_, new_n_n682_, new_n_n1683_, new_n_n651_, new_n_n643_,
    new_n_n634_, new_n_n626_, new_n_n1670_, new_n_n592_, new_n_n572_,
    new_n_n570_, new_n_n562_, new_n_n551_, new_n_n1658_, new_n_n516_,
    new_n_n507_, new_n_n496_, new_n_n1648_, new_n_n485_, new_n_n476_,
    new_n_n1646_, new_n_n457_, new_n_n1639_, new_n_n424_, new_n_n414_,
    new_n_n407_, new_n_n403_, new_n_n395_, new_n_n383_, new_n_n375_,
    new_n_n349_, new_n_n341_, new_n_n1618_, new_n_n324_, new_n_n1615_,
    new_n_n311_, new_n_n299_, new_n_n291_, new_n_n266_, new_n_n261_,
    new_n_n253_, new_n_n241_, new_n_n232_, new_n_n228_, new_n_n207_,
    new_n_n198_, new_n_n1605_, new_n_n173_, new_n_n1604_, new_n_n160_,
    new_n_n148_, new_n_n140_, new_n_n115_, new_n_n106_, new_n_n2_,
    new_n_n1594_, new_n_n2470_, new_n_n2465_, new_n_n2432_, new_n_n2424_,
    new_n_n2419_, new_n_n2410_, new_n_n2405_, new_n_n2397_, new_n_n1565_,
    new_n_n2378_, new_n_n1550_, new_n_n2369_, new_nb14_, new_n_n1538_,
    new_n_n2353_, new_nb13_, new_n_n2344_, new_n_n1515_, new_n_n1512_,
    new_n_n2322_, new_n_n1504_, new_n_n2314_, new_n_n1495_, new_n_n1491_,
    new_n_n2284_, new_n_n2280_, new_n_n2276_, new_n_n2267_, new_n_n2237_,
    new_n_n2009_, new_n_n1174_, new_n_n1980_, new_n_n1974_, new_n_n1133_,
    new_n_n1966_, new_n_n1122_, new_n_n1105_, new_n_n1943_, new_n_n1940_,
    new_n_n1090_, new_n_n1930_, new_n_n1080_, new_n_n1924_, new_n_n1918_,
    new_n_n1912_, new_n_n1058_, new_n_n1057_, new_n_n1051_, new_n_n1048_,
    new_n_n1888_, new_n_n1038_, new_n_n1032_, new_n_n1023_, new_n_n1016_,
    new_n_n1861_, new_n_n1006_, new_n_n998_, new_n_n1853_, new_n_n987_,
    new_n_n1823_, new_n_n1819_, new_n_n949_, new_n_n815_, new_n_n804_,
    new_n_n1710_, new_n_n790_, new_n_n746_, new_n_n729_, new_n_n722_,
    new_n_n716_, new_n_n706_, new_n_n666_, new_n_n657_, new_n_n650_,
    new_n_n1677_, new_n_n636_, new_n_n627_, new_n_n1669_, new_n_n583_,
    new_n_n573_, new_n_n569_, new_n_n559_, new_n_n1659_, new_n_n543_,
    new_n_n515_, new_n_n505_, new_n_n499_, new_n_n490_, new_n_n484_,
    new_n_n473_, new_n_n467_, new_n_n458_, new_n_n443_, new_n_n1638_,
    new_n_n422_, new_n_n417_, new_n_n408_, new_n_n402_, new_n_n1629_,
    new_n_n386_, new_n_n376_, new_n_n364_, new_n_n355_, new_n_n348_,
    new_n_n338_, new_n_n333_, new_n_n325_, new_n_n319_, new_n_n308_,
    new_n_n302_, new_n_n292_, new_n_n277_, new_n_n267_, new_n_n260_,
    new_n_n250_, new_n_n1609_, new_n_n233_, new_n_n227_, new_n_n217_,
    new_n_n199_, new_n_n184_, new_n_n174_, new_n_n168_, new_n_n157_,
    new_n_n151_, new_n_n141_, new_n_n134_, new_n_n124_, new_n_n3_,
    new_n_n1596_, new_n_n1593_, new_n_n2471_, new_n_n2464_, new_n_n1578_,
    new_n_n2425_, new_n_n2418_, new_n_n2411_, new_n_n2404_, new_n_n1567_,
    new_n_n2391_, new_n_n1559_, new_n_n2377_, new_n_n1551_, new_n_n2368_,
    new_n_n2363_, new_n_n2360_, new_n_n2354_, new_n_n2349_, new_n_n2345_,
    new_n_n2339_, new_n_n2332_, new_n_n2327_, new_n_n1507_, new_n_n1503_,
    new_n_n1498_, new_n_n2309_, new_n_n2304_, new_n_n1469_, new_nb0_,
    new_n_n2277_, new_n_n2272_, new_n_n1422_, new_n_n2008_, new_n_n1175_,
    new_no9_, new_n_n1138_, new_n_n1969_, new_n_n1965_, new_n_n1123_,
    new_n_n1104_, new_n_n1944_, new_n_n1939_, new_n_n1934_, new_n_n1086_,
    new_n_n1081_, new_n_n1923_, new_n_n1072_, new_n_n1911_, new_n_n1059_,
    new_n_n1056_, new_n_n1897_, new_n_n1047_, new_n_n1043_, new_n_n1885_,
    new_n_n1033_, new_n_n1029_, new_n_n1866_, new_n_n1862_, new_n_n1005_,
    new_n_n1856_, new_n_n1852_, new_n_n988_, new_n_n964_, new_n_n959_,
    new_n_n1814_, new_n_n814_, new_n_n805_, new_n_n799_, new_n_n791_,
    new_n_n1700_, new_n_n728_, new_n_n723_, new_n_n715_, new_n_n707_,
    new_n_n665_, new_n_n658_, new_n_n649_, new_n_n1678_, new_n_n635_,
    new_n_n1674_, new_n_n590_, new_n_n582_, new_n_n574_, new_n_n568_,
    new_n_n560_, new_n_n553_, new_n_n544_, new_n_n514_, new_n_n1652_,
    new_n_n498_, new_n_n491_, new_n_n483_, new_n_n474_, new_n_n466_,
    new_n_n459_, new_n_n435_, new_n_n1637_, new_n_n1636_, new_n_n416_,
    new_n_n1632_, new_n_n401_, new_n_n393_, new_n_n385_, new_n_n1628_,
    new_n_n363_, new_n_n356_, new_n_n347_, new_n_n339_, new_n_n332_,
    new_n_n326_, new_n_n318_, new_n_n309_, new_n_n301_, new_n_n293_,
    new_n_n276_, new_n_n268_, new_n_n259_, new_n_n251_, new_n_n243_,
    new_n_n234_, new_n_n226_, new_n_n1607_, new_n_n209_, new_n_n183_,
    new_n_n175_, new_n_n167_, new_n_n158_, new_n_n150_, new_n_n142_,
    new_n_n133_, new_n_n125_, new_n_n4_, new_n_n2482_, new_n_n1592_,
    new_n_n2466_, new_n_n2393_, new_n_n1372_, new_n_n1366_, new_n_n2174_,
    new_n_n1323_, new_n_n1317_, new_n_n2132_, new_n_n2126_, new_n_n1303_,
    new_n_n1297_, new_n_n2093_, new_n_n1271_, new_n_n1265_, new_n_n1258_,
    new_n_n2077_, new_n_n1243_, new_no12_, new_n_n2065_, new_n_n1226_,
    new_n_n1211_, new_n_n2037_, new_n_n1199_, new_n_n1194_, new_n_n1188_,
    new_n_n1182_, new_n_n1179_, new_ne10_, new_n_n1148_, new_n_n1977_,
    new_n_n1137_, new_n_n1130_, new_n_n1962_, new_no7_, new_n_n1919_,
    new_n_n92_, new_n_n82_, new_n_n71_, new_n_n60_, new_n_n49_,
    new_n_n2481_, new_n_n2475_, new_n_n1589_, new_n_n2392_, new_n_n1371_,
    new_n_n2180_, new_n_n2171_, new_n_n1322_, new_n_n1318_, new_n_n2131_,
    new_n_n1306_, new_n_n1302_, new_n_n2114_, new_n_n2092_, new_ne13_,
    new_n_n1264_, new_n_n2081_, new_n_n1250_, new_n_n2074_, new_n_n1236_,
    new_n_n1231_, new_n_n2055_, new_n_n2042_, new_n_n1206_, new_n_n2033_,
    new_n_n2029_, new_n_n2023_, new_n_n1183_, new_n_n2010_, new_n_n1176_,
    new_n_n1985_, new_n_n1976_, new_n_n1971_, new_n_n1129_, new_n_n1124_,
    new_n_n1077_, new_n_n1920_, new_n_n93_, new_n_n81_, new_n_n72_,
    new_n_n59_, new_n_n50_, new_n_n2480_, new_n_n2473_, new_n_n2468_,
    new_n_n2408_, new_n_n2400_, new_n_n2185_, new_n_n2181_, new_n_n2164_,
    new_n_n1324_, new_n_n2137_, new_n_n1310_, new_n_n2124_, new_n_n2119_,
    new_n_n1298_, new_n_n1272_, new_n_n2084_, new_n_n2080_, new_n_n1252_,
    new_n_n1244_, new_n_n1235_, new_n_n1227_, new_n_n2056_, new_n_n1210_,
    new_n_n2036_, new_n_n2034_, new_n_n2030_, new_n_n1187_, new_n_n2017_,
    new_n_n2012_, new_n_n1177_, new_n_n1157_, new_n_n1141_, new_n_n1136_,
    new_n_n1131_, new_n_n1125_, new_n_n1088_, new_n_n1083_, new_n_n94_,
    new_n_n80_, new_n_n69_, new_n_n62_, new_n_n51_, new_n_n1595_,
    new_n_n2474_, new_n_n2467_, new_n_n2407_, new_n_n1568_, new_n_n1373_,
    new_n_n2182_, new_n_n2160_, new_ne15_, new_n_n2138_, new_n_n2130_,
    new_n_n2125_, new_n_n2118_, new_n_n1299_, new_n_n1277_, new_n_n2083_,
    new_n_n1257_, new_n_n1251_, new_n_n1245_, new_n_n2064_, new_n_n2059_,
    new_n_n1220_, new_n_n1209_, new_n_n1205_, new_n_n1200_, new_n_n1195_,
    new_n_n1186_, new_n_n2018_, new_n_n2011_, new_n_n2004_, new_n_n1164_,
    new_n_n1140_, new_n_n1970_, new_n_n1967_, new_n_n1963_, new_n_n1932_,
    new_n_n1927_, new_n_n95_, new_n_n79_, new_n_n70_, new_n_n61_,
    new_n_n52_, new_n_n0_, new_n_n2423_, new_n_n2415_, new_n_n1419_,
    new_n_n2229_, new_n_n1410_, new_n_n1375_, new_n_n2183_, new_n_n2156_,
    new_n_n2141_, new_n_n1319_, new_n_n2110_, new_n_n2104_, new_n_n2100_,
    new_n_n1278_, new_n_n1263_, new_n_n1255_, new_n_n1248_, new_n_n2071_,
    new_n_n1232_, new_n_n2060_, new_n_n2057_, new_n_n2041_, new_n_n1204_,
    new_n_n2032_, new_n_n2026_, new_n_n1190_, new_n_n1185_, new_n_n2014_,
    new_n_n2005_, new_n_n1163_, new_n_n1989_, new_n_n1151_, new_n_n1145_,
    new_n_n1126_, new_n_n1942_, new_n_n1937_, new_n_n1775_, new_n_n903_,
    new_n_n803_, new_n_n1709_, new_n_n1694_, new_n_n1599_, new_n_n42_,
    new_n_n31_, new_n_n20_, new_n_n9_, new_n_n1590_, new_n_n1575_,
    new_n_n2416_, new_n_n1467_, new_n_n1420_, new_n_n2228_, new_n_n2222_,
    new_n_n1374_, new_n_n1367_, new_n_n2150_, new_n_n1325_, new_no15_,
    new_n_n1294_, new_n_n1290_, new_n_n2099_, new_n_n2094_, new_n_n2082_,
    new_n_n1256_, new_n_n1241_, new_n_n2070_, new_n_n1233_, new_n_n1228_,
    new_n_n1221_, new_n_n2040_, new_n_n2035_, new_n_n2031_, new_n_n1193_,
    new_n_n2025_, new_n_n2020_, new_n_n2013_, new_n_n2006_, new_n_n1162_,
    new_n_n1990_, new_n_n1983_, new_n_n1146_, new_n_n1132_, new_n_n1098_,
    new_n_n1093_, new_n_n1774_, new_n_n904_, new_n_n802_, new_n_n796_,
    new_n_n720_, new_n_n96_, new_n_n41_, new_n_n32_, new_n_n19_,
    new_n_n10_, new_n_n2476_, new_n_n2438_, new_n_n2430_, new_n_n1461_,
    new_nb5_, new_n_n1414_, new_n_n2223_, new_nb10_, new_n_n1368_,
    new_n_n1331_, new_n_n1293_, new_n_n1288_, new_n_n2101_, new_n_n2095_,
    new_n_n1262_, new_n_n1249_, new_n_n2073_, new_n_n1238_, new_n_n2066_,
    new_n_n2062_, new_n_n1222_, new_n_n1208_, new_ne11_, new_no11_,
    new_n_n2027_, new_n_n2024_, new_n_n1184_, new_n_n1180_, new_n_n1178_,
    new_n_n1993_, new_n_n1156_, new_n_n1984_, new_ne9_, new_n_n1972_,
    new_n_n1952_, new_n_n1947_, new_n_n961_, new_n_n909_, new_ne1_,
    new_n_n820_, new_n_n812_, new_n_n1698_, new_n_n40_, new_n_n29_,
    new_n_n22_, new_n_n11_, new_n_n2483_, new_n_n1580_, new_n_n2431_,
    new_n_n1456_, new_n_n2233_, new_n_n2230_, new_n_n2224_, new_n_n2186_,
    new_n_n1369_, new_n_n2142_, new_n_n1292_, new_n_n1289_, new_n_n1283_,
    new_n_n2096_, new_n_n2079_, new_n_n2076_, new_n_n1242_, new_n_n1237_,
    new_n_n2067_, new_n_n2061_, new_n_n1223_, new_n_n2039_, new_n_n1203_,
    new_n_n1198_, new_n_n2028_, new_n_n1189_, new_n_n2019_, new_n_n2015_,
    new_n_n2007_, new_n_n1161_, new_n_n1988_, new_n_n1152_, new_n_n1147_,
    new_n_n1142_, new_n_n1108_, new_n_n1103_, new_n_n956_, new_n_n1776_,
    new_n_n905_, new_n_n1715_, new_n_n813_, new_n_n736_, new_n_n39_,
    new_n_n30_, new_n_n21_, new_n_n12_, new_n_n1585_, new_n_n2445_,
    new_n_n1451_, new_n_n1406_, new_n_n1400_, new_n_n1395_, new_n_n2203_,
    new_n_n1364_, new_n_n1360_, new_n_n1354_, new_n_n2162_, new_n_n1344_,
    new_n_n2151_, new_n_n1332_, new_n_n1326_, new_n_n1305_, new_n_n2116_,
    new_no14_, new_n_n2107_, new_n_n1285_, new_n_n1279_, new_n_n1273_,
    new_n_n2069_, new_n_n1229_, new_n_n1224_, new_n_n1217_, new_n_n2045_,
    new_n_n2002_, new_n_n1997_, new_n_n1120_, new_no8_, new_n_n950_,
    new_n_n898_, new_n_n893_, new_n_n888_, new_n_n881_, new_n_n1720_,
    new_n_n827_, new_n_n745_, new_n_n68_, new_n_n57_, new_n_n46_,
    new_n_n35_, new_n_n24_, new_n_n13_, new_n_n2453_, new_n_n2446_,
    new_n_n2261_, new_n_n2219_, new_n_n1401_, new_n_n1394_, new_n_n1390_,
    new_n_n2178_, new_n_n2173_, new_n_n1353_, new_n_n1349_, new_n_n1343_,
    new_n_n2152_, new_n_n2147_, new_n_n2143_, new_n_n1304_, new_n_n2117_,
    new_n_n1295_, new_n_n1291_, new_n_n1284_, new_n_n1280_, new_n_n1267_,
    new_n_n1240_, new_n_n2063_, new_n_n2058_, new_n_n1216_, new_n_n1212_,
    new_no10_, new_n_n1167_, new_n_n1119_, new_n_n1114_, new_n_n1806_,
    new_n_n897_, new_n_n1764_, new_n_n1757_, new_n_n882_, new_n_n835_,
    new_n_n828_, new_n_n754_, new_n_n67_, new_n_n58_, new_n_n45_,
    new_n_n36_, new_n_n23_, new_n_n14_, new_n_n2460_, new_n_n1443_,
    new_n_n1405_, new_n_n1399_, new_n_n1396_, new_n_n2204_, new_n_n2177_,
    new_n_n2172_, new_n_n2169_, new_n_n1350_, new_n_n1342_, new_n_n1337_,
    new_n_n2149_, new_n_n1327_, new_n_n2134_, new_n_n2128_, new_n_n2112_,
    new_n_n2105_, new_n_n1287_, new_n_n1281_, new_n_n2090_, new_no13_,
    new_n_n1239_, new_n_n1234_, new_n_n1225_, new_n_n2051_, new_n_n1213_,
    new_n_n1173_, new_n_n1998_, new_n_n940_, new_n_n1768_, new_n_n891_,
    new_n_n1759_, new_n_n1754_, new_n_n848_, new_n_n841_, new_n_n763_,
    new_n_n88_, new_n_n77_, new_n_n44_, new_n_n33_, new_n_n26_, new_n_n15_,
    new_n_n2461_, new_n_n1438_, new_n_n1404_, new_n_n2214_, new_n_n2209_,
    new_n_n1391_, new_n_n2176_, new_n_n1359_, new_n_n2168_, new_n_n1351_,
    new_n_n1341_, new_n_n1338_, new_n_n2148_, new_n_n1328_, new_n_n1314_,
    new_n_n2129_, new_n_n2111_, new_n_n2106_, new_n_n1286_, new_n_n2097_,
    new_n_n2089_, new_n_n2087_, new_n_n2072_, new_n_n2068_, new_n_n1230_,
    new_n_n1218_, new_n_n2046_, new_n_n1172_, new_n_n1999_, new_ne2_,
    new_no1_, new_n_n892_, new_n_n1758_, new_n_n1755_, new_n_n847_,
    new_n_n1724_, new_n_n1706_, new_n_n87_, new_n_n78_, new_n_n43_,
    new_n_n34_, new_n_n25_, new_n_n16_, new_n_n2246_, new_n_n2199_,
    new_n_n2194_, new_n_n1377_, new_n_n2175_, new_n_n1357_, new_n_n2166_,
    new_n_n1347_, new_n_n2158_, new_n_n2153_, new_n_n1334_, new_n_n2144_,
    new_n_n1320_, new_n_n1315_, new_n_n1313_, new_n_n2127_, new_n_n2121_,
    new_ne14_, new_n_n2103_, new_n_n1282_, new_n_n1275_, new_n_n1268_,
    new_n_n1261_, new_n_n1253_, new_n_n1246_, new_n_n2052_, new_n_n2047_,
    new_n_n1168_, new_n_n1793_, new_n_n876_, new_n_n1747_, new_n_n863_,
    new_n_n1736_, new_n_n860_, new_n_n855_, new_n_n779_, new_n_n89_,
    new_n_n86_, new_n_n75_, new_n_n64_, new_n_n53_, new_n_n28_, new_n_n17_,
    new_n_n2243_, new_nb11_, new_n_n2195_, new_n_n1376_, new_n_n1363_,
    new_n_n1358_, new_n_n2165_, new_n_n1348_, new_n_n1346_, new_n_n2154_,
    new_n_n1333_, new_n_n1329_, new_n_n2139_, new_n_n2135_, new_n_n1312_,
    new_n_n1309_, new_n_n2120_, new_n_n1300_, new_n_n2102_, new_n_n2098_,
    new_n_n1274_, new_n_n1269_, new_n_n2086_, new_n_n2078_, new_n_n2075_,
    new_n_n1219_, new_n_n1214_, new_n_n2003_, new_n_n1788_, new_n_n875_,
    new_n_n1748_, new_n_n862_, new_n_n1737_, new_n_n1735_, new_n_n1730_,
    new_n_n788_, new_n_n1598_, new_n_n85_, new_n_n76_, new_n_n63_,
    new_n_n54_, new_n_n27_, new_n_n18_, new_n_n2238_, new_n_n2198_,
    new_n_n1381_, new_n_n2188_, new_n_n1370_, new_n_n1362_, new_n_n1355_,
    new_n_n2167_, new_n_n2161_, new_n_n1345_, new_n_n1339_, new_n_n1336_,
    new_n_n2145_, new_n_n2140_, new_n_n2136_, new_n_n2133_, new_n_n1307_,
    new_n_n2123_, new_n_n1301_, new_n_n1296_, new_n_n2108_, new_n_n1276_,
    new_n_n2088_, new_n_n2085_, new_n_n1259_, new_n_n1247_, new_n_n2054_,
    new_n_n1215_, new_n_n918_, new_n_n1751_, new_n_n868_, new_n_n864_,
    new_n_n1738_, new_n_n90_, new_n_n84_, new_n_n73_, new_n_n66_,
    new_n_n55_, new_n_n48_, new_n_n37_, new_n_n1386_, new_n_n2193_,
    new_n_n1378_, new_n_n1365_, new_n_n1361_, new_n_n1356_, new_n_n1352_,
    new_nb8_, new_n_n2157_, new_n_n1340_, new_n_n1335_, new_n_n2146_,
    new_n_n1321_, new_n_n1316_, new_n_n1311_, new_n_n1308_, new_n_n2122_,
    new_n_n2115_, new_n_n2113_, new_n_n2109_, new_n_n2091_, new_n_n1270_,
    new_n_n1266_, new_n_n1260_, new_n_n1254_, new_n_n2053_, new_n_n2048_,
    new_n_n913_, new_n_n874_, new_n_n869_, new_n_n1744_, new_n_n1739_,
    new_n_n91_, new_n_n83_, new_n_n74_, new_n_n65_, new_n_n56_, new_n_n47_,
    new_n_n38_;
  assign po12 = new_no12_;
  assign new_nina0_ = pina0;
  assign new_ninb1_ = pinb1;
  assign new_ninc2_ = pinc2;
  assign new_nind3_ = pind3;
  assign po11 = new_no11_;
  assign new_nina1_ = pina1;
  assign new_ninb0_ = pinb0;
  assign new_ninc3_ = pinc3;
  assign new_nind2_ = pind2;
  assign new_nmusel1_ = pmusel1;
  assign po14 = new_no14_;
  assign new_ninc4_ = pinc4;
  assign new_nind5_ = pind5;
  assign new_nmusel2_ = pmusel2;
  assign po13 = new_no13_;
  assign new_ninc5_ = pinc5;
  assign new_nind4_ = pind4;
  assign new_nmusel3_ = pmusel3;
  assign new_nina4_ = pina4;
  assign new_ninb5_ = pinb5;
  assign po15 = new_no15_;
  assign new_nina5_ = pina5;
  assign new_ninb4_ = pinb4;
  assign po9 = new_no9_;
  assign new_nina2_ = pina2;
  assign new_ninb3_ = pinb3;
  assign new_ninc0_ = pinc0;
  assign new_nind1_ = pind1;
  assign po8 = new_no8_;
  assign new_nina3_ = pina3;
  assign new_ninb2_ = pinb2;
  assign new_ninc1_ = pinc1;
  assign new_nind0_ = pind0;
  assign po7 = new_no7_;
  assign po6 = new_no6_;
  assign new_nind15_ = pind15;
  assign po5 = new_no5_;
  assign new_ninc15_ = pinc15;
  assign new_nind14_ = pind14;
  assign po4 = new_no4_;
  assign new_ninb15_ = pinb15;
  assign new_ninc14_ = pinc14;
  assign new_nind13_ = pind13;
  assign po3 = new_no3_;
  assign new_nopsel3_ = popsel3;
  assign po2 = new_no2_;
  assign po1 = new_no1_;
  assign new_nopsel1_ = popsel1;
  assign po0 = new_no0_;
  assign new_nopsel2_ = popsel2;
  assign new_nina11_ = pina11;
  assign new_ninb10_ = pinb10;
  assign new_nina10_ = pina10;
  assign new_nopsel0_ = popsel0;
  assign new_nina15_ = pina15;
  assign new_ninb14_ = pinb14;
  assign new_ninc13_ = pinc13;
  assign new_nind12_ = pind12;
  assign new_nina14_ = pina14;
  assign new_ninb13_ = pinb13;
  assign new_ninc12_ = pinc12;
  assign new_nind11_ = pind11;
  assign new_nina13_ = pina13;
  assign new_ninb12_ = pinb12;
  assign new_ninc11_ = pinc11;
  assign new_nind10_ = pind10;
  assign new_nina12_ = pina12;
  assign new_ninb11_ = pinb11;
  assign new_ninc10_ = pinc10;
  assign new_nina8_ = pina8;
  assign new_ninb9_ = pinb9;
  assign new_nina9_ = pina9;
  assign new_ninb8_ = pinb8;
  assign new_nina6_ = pina6;
  assign new_ninb7_ = pinb7;
  assign new_nina7_ = pina7;
  assign new_ninb6_ = pinb6;
  assign new_nsh0_ = psh0;
  assign new_ninc6_ = pinc6;
  assign new_nind7_ = pind7;
  assign new_nmusel4_ = pmusel4;
  assign new_nsh1_ = psh1;
  assign new_ninc7_ = pinc7;
  assign new_nind6_ = pind6;
  assign new_nsh2_ = psh2;
  assign po10 = new_no10_;
  assign new_ninc8_ = pinc8;
  assign new_nind9_ = pind9;
  assign new_ninc9_ = pinc9;
  assign new_nind8_ = pind8;
  assign new_n_n2456_ = new_n_n24_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n1583_ = new_n_n31_ & new_n_n840_;
  assign new_n_n2439_ = new_n_n1714_ | new_n_n815_ | new_n_n282_;
  assign new_n_n2385_ = new_n_n1724_ | new_n_n1635_;
  assign new_n_n2380_ = new_n_n89_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2372_ = new_n_n1549_ | new_n_n1551_ | new_n_n1550_ | new_n_n893_;
  assign new_n_n1546_ = new_n_n107_ & new_n_n108_;
  assign new_n_n1542_ = new_n_n2159_ & new_nb14_;
  assign new_n_n1536_ = new_n_n1714_ & new_n_n119_;
  assign new_n_n1517_ = new_n_n142_ & new_n_n1715_;
  assign new_n_n2329_ = new_n_n848_ & new_n_n1730_ & new_n_n853_;
  assign new_n_n1508_ = new_n_n1714_ & new_n_n151_;
  assign new_n_n2317_ = new_n_n159_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2312_ = new_n_n1715_ | new_n_n820_ | new_n_n751_;
  assign new_n_n1493_ = new_n_n170_ & new_n_n1714_;
  assign new_n_n1486_ = new_n_n770_ & new_n_n728_;
  assign new_n_n2297_ = new_n_n1480_ | new_n_n819_;
  assign new_n_n2291_ = new_n_n1475_ | new_n_n1476_;
  assign new_n_n1460_ = new_n_n845_ & new_n_n801_;
  assign new_n_n2271_ = new_n_n728_ | new_n_n1699_;
  assign new_n_n2265_ = new_n_n1715_ | new_n_n820_ | new_n_n580_;
  assign new_n_n1446_ = new_n_n219_ & new_n_n1714_;
  assign new_n_n2255_ = new_n_n225_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2247_ = new_n_n1434_ | new_n_n1436_ | new_n_n1435_ | new_n_n893_;
  assign new_n_n1430_ = new_n_n1678_ & new_n_n598_;
  assign new_n_n1424_ = new_n_n1714_ & new_n_n239_;
  assign new_n_n1398_ = new_n_n269_ & new_n_n642_;
  assign new_n_n2208_ = new_n_n275_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2200_ = new_n_n1387_ | new_n_n1389_ | new_n_n1388_ | new_n_n893_;
  assign new_n_n1383_ = new_n_n295_ & new_n_n1715_;
  assign new_n_n2190_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n293_;
  assign new_n_n1330_ = new_n_n344_ & new_n_n338_;
  assign new_n_n1956_ = new_n_n1114_ | new_n_n1115_;
  assign new_n_n1953_ = new_n_n1665_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1064_ = new_n_n631_ & new_n_n1721_;
  assign new_n_n1907_ = new_n_n1058_ | new_n_n1059_;
  assign new_n_n1900_ = new_n_n645_ | new_n_n1679_;
  assign new_n_n1896_ = new_n_n653_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n1891_ = new_n_n1719_ | new_n_n1681_;
  assign new_n_n1868_ = new_n_n1685_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1011_ = new_n_n665_ & new_n_n1720_;
  assign new_n_n1858_ = new_n_n1003_ | new_n_n1004_;
  assign new_n_n1855_ = new_n_n994_ | new_n_n913_ | new_n_n995_ | new_n_n996_;
  assign new_n_n990_ = new_n_n708_ & new_n_n1730_;
  assign new_n_n985_ = new_n_n786_ & new_n_n1719_;
  assign new_n_n1841_ = new_n_n977_ | new_n_n978_;
  assign new_n_n1836_ = new_n_n1724_ | new_n_n724_;
  assign new_n_n960_ = new_n_n751_ & new_n_n1714_;
  assign new_n_n955_ = new_n_n833_ & new_n_n757_;
  assign new_n_n1809_ = new_n_n764_ | new_n_n765_;
  assign new_n_n943_ = new_n_n768_ & new_n_n769_;
  assign new_n_n937_ = new_n_n1727_ & new_n_n734_;
  assign new_n_n1795_ = new_n_n777_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n1790_ = new_n_n1719_ | new_n_n1708_;
  assign new_n_n1785_ = new_n_n883_ | new_n_n879_ | new_n_n918_ | new_n_n919_;
  assign new_n_n914_ = new_n_n853_ & new_n_n1710_;
  assign new_n_n890_ = new_n_n817_ & new_n_n818_;
  assign new_n_n886_ = new_n_n831_ & new_n_n826_;
  assign new_n_n879_ = new_n_n833_ & new_n_n1720_;
  assign new_n_n871_ = new_n_n841_ & new_n_n1725_;
  assign new_ne0_ = new_n_n864_ | new_n_n865_;
  assign new_n_n1740_ = new_n_n1638_ & new_n_n2337_;
  assign new_n_n858_ = ~new_n_n1726_;
  assign new_n_n851_ = ~new_ne0_;
  assign new_n_n1725_ = ~new_n_n1752_;
  assign new_n_n838_ = ~new_n_n1753_;
  assign new_n_n1718_ = ~new_n_n1760_;
  assign new_n_n1716_ = ~new_nmusel4_;
  assign new_n_n785_ = ~new_n_n1790_;
  assign new_n_n775_ = ~new_n_n1704_;
  assign new_n_n767_ = ~new_n_n1806_;
  assign new_n_n758_ = ~new_n_n1650_;
  assign new_n_n748_ = ~new_n_n1822_;
  assign new_n_n737_ = ~new_n_n1798_;
  assign new_n_n1699_ = ~new_n_n2322_;
  assign new_n_n1692_ = ~new_n_n2442_;
  assign new_n_n696_ = ~new_n_n1688_;
  assign new_n_n686_ = ~new_n_n1868_;
  assign new_n_n676_ = ~new_n_n1873_;
  assign new_n_n668_ = ~new_n_n1883_;
  assign new_n_n1680_ = ~new_nind5_;
  assign new_n_n648_ = ~new_n_n1902_;
  assign new_n_n640_ = ~new_n_n1876_;
  assign new_n_n622_ = ~new_n_n1924_;
  assign new_n_n611_ = ~new_n_n1928_;
  assign new_n_n601_ = ~new_n_n2277_;
  assign new_n_n594_ = ~new_n_n1942_;
  assign new_n_n585_ = ~new_n_n1950_;
  assign new_n_n575_ = ~new_n_n1664_;
  assign new_n_n567_ = ~new_n_n1964_;
  assign new_n_n1660_ = ~new_n_n1974_;
  assign new_n_n548_ = ~new_n_n1979_;
  assign new_n_n540_ = ~new_n_n1986_;
  assign new_n_n531_ = ~new_n_n1997_;
  assign new_n_n521_ = ~new_n_n1652_;
  assign new_n_n510_ = ~new_n_n1618_;
  assign new_n_n501_ = ~new_n_n2429_;
  assign new_n_n492_ = ~new_n_n2028_;
  assign new_n_n482_ = ~new_n_n1646_;
  assign new_n_n471_ = ~new_n_n1212_;
  assign new_n_n462_ = ~new_n_n2050_;
  assign new_n_n452_ = ~new_n_n2059_;
  assign new_n_n442_ = ~new_n_n2075_;
  assign new_n_n434_ = ~new_n_n351_;
  assign new_n_n427_ = ~new_n_n2082_;
  assign new_n_n419_ = ~new_n_n2086_;
  assign new_n_n1633_ = ~new_n_n2343_;
  assign new_n_n400_ = ~new_n_n2107_;
  assign new_n_n391_ = ~new_ninb13_;
  assign new_n_n380_ = ~new_n_n2116_;
  assign new_n_n372_ = ~new_n_n2092_;
  assign new_n_n354_ = ~new_n_n2139_;
  assign new_n_n344_ = ~new_n_n1741_;
  assign new_n_n1620_ = ~new_n_n2198_;
  assign new_n_n327_ = ~new_nb8_;
  assign new_n_n317_ = ~new_n_n2168_;
  assign new_n_n1614_ = ~new_ninc9_;
  assign new_n_n296_ = ~new_n_n2189_;
  assign new_n_n286_ = ~new_n_n2202_;
  assign new_n_n256_ = ~new_n_n2225_;
  assign new_n_n245_ = ~new_nina5_;
  assign new_n_n235_ = ~new_n_n2246_;
  assign new_n_n225_ = ~new_n_n2256_;
  assign new_n_n215_ = ~new_n_n2264_;
  assign new_n_n204_ = ~new_n_n2275_;
  assign new_n_n194_ = ~new_n_n2284_;
  assign new_n_n153_ = ~new_n_n2323_;
  assign new_n_n1602_ = ~new_ninc12_;
  assign new_n_n132_ = ~new_n_n2345_;
  assign new_n_n122_ = ~new_n_n2354_;
  assign new_n_n112_ = ~new_n_n2364_;
  assign new_n_n101_ = ~new_n_n2374_;
  assign new_n_n1586_ = new_n_n23_ & new_n_n1714_;
  assign new_n_n2447_ = new_n_n1610_ | new_n_n1715_;
  assign new_n_n2440_ = new_n_n1612_ | new_n_n1715_;
  assign new_n_n1561_ = new_n_n83_ & new_n_n84_;
  assign new_n_n2379_ = new_n_n815_ | new_n_n1713_ | new_n_n1598_;
  assign new_n_n2373_ = new_n_n96_ & new_n_n815_;
  assign new_n_n2367_ = new_n_n1600_ | new_n_n1716_;
  assign new_n_n2362_ = new_n_n1541_ | new_n_n1542_;
  assign new_n_n1532_ = new_n_n129_ & new_n_n124_;
  assign new_n_n1518_ = new_n_n815_ & new_n_n1602_;
  assign new_n_n2328_ = new_n_n1512_ | new_n_n849_;
  assign new_n_n2323_ = new_n_n1507_ | new_n_n1508_;
  assign new_nb3_ = new_n_n160_ & new_n_n161_;
  assign new_n_n2313_ = new_n_n815_ | new_n_n1713_ | new_n_n1701_;
  assign new_n_n1492_ = new_n_n170_ & new_n_n171_;
  assign new_n_n1487_ = new_n_n770_ & new_n_n1699_;
  assign new_n_n1480_ = new_n_n179_ & new_n_n180_;
  assign new_nb1_ = new_n_n186_ & new_n_n187_;
  assign new_n_n1466_ = new_n_n196_ & new_n_n197_;
  assign new_n_n2270_ = new_n_n1455_ | new_n_n207_;
  assign new_n_n2266_ = new_n_n815_ | new_n_n1713_ | new_n_n1665_;
  assign new_n_n1445_ = new_n_n219_ & new_n_n220_;
  assign new_n_n1440_ = new_n_n232_ & new_n_n1608_;
  assign new_n_n1436_ = new_n_n79_ & new_n_n233_;
  assign new_n_n1431_ = new_n_n1678_ & new_n_n1670_;
  assign new_n_n1423_ = new_n_n1714_ & new_n_n240_;
  assign new_n_n2213_ = new_n_n1678_ & new_n_n642_;
  assign new_n_n1393_ = new_n_n282_ & new_n_n1612_;
  assign new_n_n1389_ = new_n_n79_ & new_n_n283_;
  assign new_n_n1384_ = new_n_n815_ & new_n_n1613_;
  assign new_n_n2189_ = new_n_n294_ & new_n_n815_;
  assign new_ng3_ = new_n_n1333_ | new_n_n1335_ | new_n_n1334_ | new_n_n1336_;
  assign new_n_n1115_ = new_n_n574_ & new_n_n351_;
  assign new_n_n1109_ = new_n_n580_ & new_n_n581_;
  assign new_n_n1913_ = new_n_n1691_ | new_n_n670_ | new_n_n1692_;
  assign new_n_n1908_ = new_n_n636_ & new_n_n351_;
  assign new_n_n1899_ = new_n_n646_ | new_n_n266_;
  assign new_n_n1050_ = new_n_n385_ & new_n_n652_;
  assign new_n_n1886_ = new_n_n1011_ | new_n_n879_ | new_n_n1038_ | new_n_n1039_;
  assign new_n_n1867_ = new_n_n1016_ | new_n_n686_;
  assign new_n_n1012_ = new_n_n665_ & new_n_n689_;
  assign new_n_n1004_ = new_n_n1689_ & new_n_n697_;
  assign new_n_n997_ = new_n_n701_ & new_n_n1692_;
  assign new_n_n1851_ = new_n_n709_ & new_n_n815_;
  assign new_n_n1846_ = new_n_n985_ | new_n_n714_;
  assign new_n_n978_ = new_n_n836_ & new_n_n719_;
  assign new_n_n973_ = new_n_n724_ & new_n_n1724_;
  assign new_n_n965_ = new_n_n743_ & new_n_n744_;
  assign new_n_n954_ = new_n_n718_ & new_n_n757_;
  assign new_n_n1810_ = new_n_n840_ | new_n_n795_ | new_n_n1722_;
  assign new_n_n1803_ = new_n_n2297_ | new_n_n1711_;
  assign new_n_n1799_ = new_n_n937_ | new_n_n772_;
  assign new_no2_ = new_n_n930_ | new_n_n778_;
  assign new_n_n926_ = new_n_n83_ & new_n_n784_;
  assign new_n_n919_ = new_n_n833_ & new_n_n789_;
  assign new_n_n1780_ = new_n_n911_ | new_n_n913_ | new_n_n912_ | new_n_n914_;
  assign new_n_n1763_ = new_n_n1713_ | new_n_n819_;
  assign new_n_n887_ = new_n_n825_ & new_n_n1719_;
  assign new_n_n878_ = new_n_n835_ & new_n_n834_;
  assign new_n_n872_ = new_n_n853_ & new_n_n1725_;
  assign new_n_n865_ = new_n_n846_ & new_n_n1727_;
  assign new_n_n1741_ = new_n_n1732_ & new_n_n857_;
  assign new_n_n1733_ = ~new_n_n2279_;
  assign new_n_n852_ = ~new_n_n1744_;
  assign new_n_n844_ = ~new_n_n1723_;
  assign new_n_n1721_ = ~new_nsh0_;
  assign new_n_n829_ = ~new_n_n1660_;
  assign new_n_n1717_ = ~new_nind0_;
  assign new_n_n784_ = ~new_n_n1793_;
  assign new_n_n776_ = ~new_ne2_;
  assign new_n_n766_ = ~new_n_n1808_;
  assign new_n_n1702_ = ~new_n_n1818_;
  assign new_n_n747_ = ~new_n_n1823_;
  assign new_n_n738_ = ~new_n_n1832_;
  assign new_n_n721_ = ~new_n_n1839_;
  assign new_n_n701_ = ~new_n_n1691_;
  assign new_n_n1687_ = ~new_n_n2220_;
  assign new_n_n1685_ = ~new_nind4_;
  assign new_n_n677_ = ~new_n_n1875_;
  assign new_n_n667_ = ~new_n_n1886_;
  assign new_n_n659_ = ~new_n_n1893_;
  assign new_n_n647_ = ~new_n_n1899_;
  assign new_n_n641_ = ~new_n_n1903_;
  assign new_n_n621_ = ~new_ninb6_;
  assign new_n_n612_ = ~new_n_n1937_;
  assign new_n_n600_ = ~new_n_n1671_;
  assign new_n_n595_ = ~new_n_n1940_;
  assign new_n_n584_ = ~new_n_n1951_;
  assign new_n_n576_ = ~new_n_n1961_;
  assign new_n_n566_ = ~new_n_n1661_;
  assign new_n_n558_ = ~new_n_n1969_;
  assign new_n_n541_ = ~new_n_n1985_;
  assign new_n_n539_ = ~new_n_n1988_;
  assign new_n_n532_ = ~new_n_n1996_;
  assign new_n_n520_ = ~new_n_n2007_;
  assign new_n_n511_ = ~new_n_n1647_;
  assign new_n_n500_ = ~new_n_n2022_;
  assign new_n_n1649_ = ~new_n_n2066_;
  assign new_n_n481_ = ~new_n_n2040_;
  assign new_n_n472_ = ~new_n_n2014_;
  assign new_n_n461_ = ~new_n_n2052_;
  assign new_n_n453_ = ~new_n_n1133_;
  assign new_n_n451_ = ~new_n_n2060_;
  assign new_n_n433_ = ~new_n_n2076_;
  assign new_n_n428_ = ~new_n_n2079_;
  assign new_n_n418_ = ~new_ninb12_;
  assign new_n_n409_ = ~new_n_n1732_;
  assign new_n_n399_ = ~new_n_n2102_;
  assign new_n_n392_ = ~new_n_n2111_;
  assign new_n_n379_ = ~new_n_n2117_;
  assign new_n_n373_ = ~new_n_n2120_;
  assign new_n_n353_ = ~new_n_n2140_;
  assign new_n_n345_ = ~new_n_n2146_;
  assign new_n_n1619_ = ~new_n_n2204_;
  assign new_n_n1616_ = ~new_n_n2043_;
  assign new_n_n316_ = ~new_n_n2169_;
  assign new_n_n307_ = ~new_n_n1614_;
  assign new_n_n295_ = ~new_nina10_;
  assign new_n_n287_ = ~new_nb11_;
  assign new_n_n265_ = ~new_n_n2219_;
  assign new_n_n244_ = ~new_n_n1609_;
  assign new_n_n236_ = ~new_n_n2249_;
  assign new_n_n224_ = ~new_nb7_;
  assign new_n_n216_ = ~new_n_n2267_;
  assign new_n_n203_ = ~new_n_n2278_;
  assign new_n_n1606_ = ~new_ninc0_;
  assign new_n_n152_ = ~new_n_n2324_;
  assign new_n_n143_ = ~new_n_n2336_;
  assign new_n_n131_ = ~new_n_n2346_;
  assign new_n_n123_ = ~new_n_n1601_;
  assign new_n_n111_ = ~new_n_n2365_;
  assign new_n_n102_ = ~new_n_n2160_;
  assign new_n_n2454_ = new_n_n1585_ | new_n_n25_;
  assign new_n_n2449_ = new_n_n840_ | new_n_n31_;
  assign new_n_n2441_ = new_n_n1692_ | new_n_n634_ | new_n_n670_ | new_n_n593_;
  assign new_n_n1560_ = new_n_n86_ & new_n_n1724_;
  assign new_n_n1556_ = new_n_n97_ & new_n_n1715_;
  assign new_n_n2374_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n95_;
  assign new_n_n2366_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n109_;
  assign new_n_n2357_ = new_n_n1536_ | new_n_n1537_;
  assign new_n_n1533_ = new_n_n129_ & new_n_n1714_;
  assign new_n_n2335_ = new_n_n143_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n1513_ = new_n_n146_ & new_n_n147_;
  assign new_n_n2324_ = new_n_n1715_ | new_n_n820_ | new_n_n710_;
  assign new_n_n2316_ = new_n_n1501_ | new_n_n1502_;
  assign new_n_n1497_ = new_n_n1714_ & new_n_n164_;
  assign new_n_n2306_ = new_n_n1492_ | new_n_n1494_ | new_n_n1493_ | new_n_n893_;
  assign new_n_n1488_ = new_n_n1706_ & new_n_n728_;
  assign new_n_n2287_ = new_n_n1715_ | new_n_n820_ | new_n_n817_;
  assign new_n_n1471_ = new_n_n1714_ & new_n_n190_;
  assign new_n_n1455_ = new_n_n208_ & new_n_n209_;
  assign new_n_n1450_ = new_n_n1714_ & new_n_n213_;
  assign new_n_n2259_ = new_n_n1445_ | new_n_n1447_ | new_n_n1446_ | new_n_n893_;
  assign new_n_n1441_ = new_n_n232_ & new_n_n1715_;
  assign new_n_n1435_ = new_n_n232_ & new_n_n1714_;
  assign new_n_n1428_ = new_n_n642_ & new_n_n598_;
  assign new_n_n2240_ = new_n_n1715_ | new_n_n820_ | new_n_n657_;
  assign new_n_n1409_ = new_n_n258_ & new_n_n1714_;
  assign new_n_n1402_ = new_n_n695_ & new_n_n675_;
  assign new_n_n1388_ = new_n_n282_ & new_n_n1714_;
  assign new_n_n2196_ = new_n_n288_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n1379_ = new_n_n291_ & new_n_n292_;
  assign new_n_n2155_ = new_n_n466_ | new_n_n1619_;
  assign new_n_n1169_ = new_n_n527_ & new_n_n1714_;
  assign new_n_n1958_ = new_n_n1724_ | new_n_n572_;
  assign new_n_n1110_ = new_n_n580_ & new_n_n1714_;
  assign new_n_n1914_ = new_n_n1064_ | new_n_n1065_;
  assign new_n_n1909_ = new_n_n1724_ | new_n_n635_;
  assign new_n_n1898_ = new_n_n1054_ | new_n_n1055_;
  assign new_n_n1892_ = new_n_n1045_ | new_n_n659_;
  assign new_n_n1887_ = new_n_n1137_ | new_n_n1015_;
  assign new_n_n1018_ = new_n_n684_ & new_n_n1714_;
  assign new_n_n1013_ = new_n_n833_ & new_n_n689_;
  assign new_n_n1003_ = new_n_n1690_ & new_n_n698_;
  assign new_n_n995_ = new_n_n703_ & new_n_n702_;
  assign new_no4_ = new_n_n990_ | new_n_n991_;
  assign new_n_n1847_ = new_n_n1719_ | new_n_n1695_;
  assign new_n_n1831_ = new_n_n2310_ | new_n_n1705_;
  assign new_n_n966_ = new_n_n743_ & new_n_n742_;
  assign new_n_n953_ = new_n_n718_ & new_n_n1720_;
  assign new_n_n948_ = new_n_n764_ & new_n_n765_;
  assign new_n_n1804_ = new_n_n943_ | new_n_n944_;
  assign new_n_n938_ = new_n_n770_ & new_n_n771_;
  assign new_n_n930_ = new_n_n779_ & new_n_n1730_;
  assign new_n_n925_ = new_n_n832_ & new_n_n1719_;
  assign new_n_n920_ = new_n_n760_ & new_n_n1720_;
  assign new_n_n915_ = new_n_n794_ & new_n_n795_;
  assign new_n_n1770_ = new_n_n899_ | new_n_n901_ | new_n_n900_ | new_n_n902_;
  assign new_n_n1767_ = new_n_n849_ | new_n_n848_;
  assign new_n_n877_ = new_n_n835_ & new_n_n1720_;
  assign new_n_n1749_ = new_n_n1724_ | new_n_n841_;
  assign new_n_n866_ = new_n_n1733_ & new_n_n1726_;
  assign new_n_n1742_ = new_n_n856_ & new_n_n1731_;
  assign new_n_n859_ = ~new_n_n1684_;
  assign new_n_n853_ = ~new_n_n1724_;
  assign new_n_n843_ = ~new_n_n1748_;
  assign new_n_n836_ = ~new_n_n1721_;
  assign new_n_n1719_ = ~new_nsh2_;
  assign new_n_n821_ = ~new_n_n1761_;
  assign new_n_n787_ = ~new_n_n1789_;
  assign new_n_n777_ = ~new_n_n1796_;
  assign new_n_n1703_ = ~new_n_n1807_;
  assign new_n_n756_ = ~new_n_n1666_;
  assign new_n_n750_ = ~new_n_n1701_;
  assign new_n_n739_ = ~new_n_n1826_;
  assign new_n_n712_ = ~new_n_n1849_;
  assign new_n_n1693_ = ~new_n_n1855_;
  assign new_n_n1688_ = ~new_n_n2226_;
  assign new_n_n685_ = ~new_n_n1870_;
  assign new_n_n1684_ = ~new_n_n2238_;
  assign new_n_n670_ = ~new_n_n2448_;
  assign new_n_n660_ = ~new_n_n1894_;
  assign new_n_n633_ = ~new_n_n1913_;
  assign new_n_n623_ = ~new_n_n1922_;
  assign new_n_n613_ = ~new_n_n1927_;
  assign new_n_n1671_ = ~new_n_n2269_;
  assign new_n_n593_ = ~new_n_n2460_;
  assign new_n_n1666_ = ~new_n_n1952_;
  assign new_n_n577_ = ~new_n_n1962_;
  assign new_n_n565_ = ~new_n_n1616_;
  assign new_n_n550_ = ~new_n_n1984_;
  assign new_n_n542_ = ~new_n_n1655_;
  assign new_n_n519_ = ~new_n_n2004_;
  assign new_n_n508_ = ~new_n_n2010_;
  assign new_n_n502_ = ~new_n_n2020_;
  assign new_n_n493_ = ~new_n_n2027_;
  assign new_n_n480_ = ~new_n_n2035_;
  assign new_n_n469_ = ~new_n_n2218_;
  assign new_n_n464_ = ~new_n_n1645_;
  assign new_n_n454_ = ~new_n_n2058_;
  assign new_n_n432_ = ~new_n_n1639_;
  assign new_n_n425_ = ~new_n_n2080_;
  assign new_n_n420_ = ~new_n_n2084_;
  assign new_n_n410_ = ~new_n_n2089_;
  assign new_n_n398_ = ~new_n_n2105_;
  assign new_n_n389_ = ~new_n_n2124_;
  assign new_n_n382_ = ~new_n_n2115_;
  assign new_n_n1626_ = ~new_n_n2362_;
  assign new_n_n352_ = ~new_ne15_;
  assign new_n_n342_ = ~new_n_n2122_;
  assign new_n_n335_ = ~new_n_n2150_;
  assign new_n_n328_ = ~new_n_n2185_;
  assign new_n_n315_ = ~new_n_n2170_;
  assign new_n_n305_ = ~new_n_n2183_;
  assign new_n_n298_ = ~new_n_n2187_;
  assign new_n_n288_ = ~new_n_n2197_;
  assign new_n_n264_ = ~new_n_n2244_;
  assign new_n_n254_ = ~new_n_n2227_;
  assign new_n_n237_ = ~new_nb6_;
  assign new_n_n223_ = ~new_n_n2261_;
  assign new_n_n213_ = ~new_n_n2266_;
  assign new_n_n206_ = ~new_n_n2274_;
  assign new_n_n195_ = ~new_n_n1606_;
  assign new_n_n171_ = ~new_n_n2307_;
  assign new_n_n161_ = ~new_n_n2320_;
  assign new_n_n130_ = ~new_n_n2348_;
  assign new_n_n120_ = ~new_n_n2357_;
  assign new_n_n114_ = ~new_n_n2366_;
  assign new_n_n103_ = ~new_n_n2161_;
  assign new_n_n2455_ = new_n_n840_ | new_n_n26_;
  assign new_n_n2448_ = new_n_n1583_ | new_n_n30_;
  assign new_n_n1581_ = new_n_n36_ & new_n_n840_;
  assign new_n_n2384_ = new_n_n1560_ | new_n_n85_;
  assign new_n_n1555_ = new_n_n97_ & new_n_n1599_;
  assign new_n_n2375_ = new_n_n1599_ | new_n_n1716_;
  assign new_n_n1541_ = new_n_n104_ & new_n_n115_;
  assign new_n_n1537_ = new_n_n1714_ & new_n_n118_;
  assign new_n_n1534_ = new_n_n79_ & new_n_n124_;
  assign new_n_n1516_ = new_n_n142_ & new_n_n1602_;
  assign new_n_n2330_ = new_n_n1729_ & new_n_n1724_ & new_n_n326_;
  assign new_n_n2325_ = new_n_n815_ | new_n_n1713_ | new_n_n1694_;
  assign new_n_n1502_ = new_n_n2159_ & new_nb3_;
  assign new_n_n2311_ = new_n_n1496_ | new_n_n1497_;
  assign new_n_n1494_ = new_n_n79_ & new_n_n171_;
  assign new_n_n1489_ = new_n_n1706_ & new_n_n1699_;
  assign new_n_n2286_ = new_n_n1470_ | new_n_n1471_;
  assign new_n_n2269_ = new_n_n1454_ | new_n_n210_;
  assign new_n_n2264_ = new_n_n1449_ | new_n_n1450_;
  assign new_n_n1447_ = new_n_n79_ & new_n_n220_;
  assign new_n_n1442_ = new_n_n815_ & new_n_n1608_;
  assign new_n_n1434_ = new_n_n232_ & new_n_n233_;
  assign new_n_n1429_ = new_n_n642_ & new_n_n1670_;
  assign new_n_n2239_ = new_n_n1423_ | new_n_n1424_;
  assign new_n_n1408_ = new_n_n258_ & new_n_n259_;
  assign new_n_n1403_ = new_n_n695_ & new_n_n1684_;
  assign new_n_n1387_ = new_n_n282_ & new_n_n283_;
  assign new_n_n1382_ = new_n_n295_ & new_n_n1613_;
  assign new_n_n2191_ = new_n_n1613_ | new_n_n1716_;
  assign new_n_n2159_ = new_n_n103_ & new_n_n1728_ & new_n_n102_;
  assign new_n_n1994_ = new_n_n1162_ | new_n_n879_ | new_n_n1163_ | new_n_n1164_;
  assign new_n_n1957_ = new_n_n573_ & new_n_n351_;
  assign new_n_n1111_ = new_n_n79_ & new_n_n581_;
  assign new_n_n1065_ = new_n_n836_ & new_n_n630_;
  assign new_n_n1060_ = new_n_n635_ & new_n_n1724_;
  assign new_no6_ = new_n_n1049_ | new_n_n654_;
  assign new_n_n1045_ = new_n_n83_ & new_n_n660_;
  assign new_n_n1040_ = new_n_n629_ & new_n_n1720_;
  assign new_n_n1017_ = new_n_n684_ & new_n_n685_;
  assign new_n_n1863_ = new_n_n1011_ | new_n_n879_ | new_n_n1012_ | new_n_n1013_;
  assign new_n_n1857_ = new_n_n999_ | new_n_n1001_ | new_n_n1000_ | new_n_n1002_;
  assign new_n_n996_ = new_n_n853_ & new_n_n702_;
  assign new_n_n991_ = new_n_n576_ & new_n_n707_;
  assign new_n_n986_ = new_n_n83_ & new_n_n713_;
  assign new_n_n1830_ = new_n_n2285_ | new_n_n1733_;
  assign new_ne3_ = new_n_n965_ | new_n_n966_;
  assign new_n_n1813_ = new_n_n1043_ | new_n_n925_;
  assign new_n_n1808_ = new_n_n948_ | new_n_n763_;
  assign new_n_n944_ = new_n_n768_ & new_n_n351_;
  assign new_n_n939_ = new_n_n1705_ & new_n_n1706_;
  assign new_n_n1794_ = new_n_n780_ & new_n_n815_;
  assign new_n_n1789_ = new_n_n925_ | new_n_n785_;
  assign new_n_n1786_ = new_n_n1014_ | new_n_n888_;
  assign new_n_n1781_ = new_n_n915_ | new_n_n793_;
  assign new_n_n902_ = new_n_n848_ & new_n_n849_;
  assign new_n_n896_ = new_n_n813_ & new_n_n1730_;
  assign new_n_n1752_ = new_n_n875_ | new_n_n876_;
  assign new_n_n870_ = new_n_n841_ & new_n_n1724_;
  assign new_n_n1745_ = new_n_n847_ & new_n_n1727_;
  assign new_n_n861_ = new_n_n855_ & new_n_n1730_;
  assign new_n_n1734_ = ~new_n_n2232_;
  assign new_n_n854_ = ~new_n_n1743_;
  assign new_n_n842_ = ~new_n_n1749_;
  assign new_n_n837_ = ~new_n_n1756_;
  assign new_n_n830_ = ~new_n_n1718_;
  assign new_n_n822_ = ~new_n_n1764_;
  assign new_n_n786_ = ~new_n_n1674_;
  assign new_n_n778_ = ~new_n_n1795_;
  assign new_n_n765_ = ~new_n_n2404_;
  assign new_n_n757_ = ~new_n_n1816_;
  assign new_n_n749_ = ~new_n_n1834_;
  assign new_n_n740_ = ~new_n_n1831_;
  assign new_n_n703_ = ~new_n_n1856_;
  assign new_n_n702_ = ~new_n_n1860_;
  assign new_n_n1689_ = ~new_n_n1859_;
  assign new_n_n684_ = ~new_ninb4_;
  assign new_n_n675_ = ~new_n_n1734_;
  assign new_n_n669_ = ~new_n_n1884_;
  assign new_n_n661_ = ~new_n_n1891_;
  assign new_n_n632_ = ~new_n_n1912_;
  assign new_n_n624_ = ~new_n_n1923_;
  assign new_n_n1673_ = ~new_nind6_;
  assign new_n_n599_ = ~new_n_n1670_;
  assign new_n_n1667_ = ~new_n_n1941_;
  assign new_n_n586_ = ~new_n_n1635_;
  assign new_n_n578_ = ~new_n_n1956_;
  assign new_n_n557_ = ~new_n_n1972_;
  assign new_n_n549_ = ~new_n_n1978_;
  assign new_n_n1656_ = ~new_n_n1991_;
  assign new_n_n518_ = ~new_n_n2009_;
  assign new_n_n509_ = ~new_n_n2008_;
  assign new_n_n1651_ = ~new_n_n2019_;
  assign new_n_n494_ = ~new_n_n1993_;
  assign new_n_n479_ = ~new_n_n2046_;
  assign new_n_n470_ = ~new_n_n2042_;
  assign new_n_n463_ = ~new_n_n2049_;
  assign new_n_n455_ = ~new_n_n2064_;
  assign new_n_n1640_ = ~new_n_n2149_;
  assign new_n_n426_ = ~new_n_n2081_;
  assign new_n_n1634_ = ~new_nind12_;
  assign new_n_n411_ = ~new_n_n2091_;
  assign new_n_n397_ = ~new_n_n2103_;
  assign new_n_n390_ = ~new_n_n1629_;
  assign new_n_n381_ = ~new_n_n2119_;
  assign new_n_n1627_ = ~new_n_n2356_;
  assign new_n_n351_ = ~new_n_n1767_;
  assign new_n_n343_ = ~new_n_n2144_;
  assign new_n_n334_ = ~new_n_n2155_;
  assign new_n_n329_ = ~new_n_n2157_;
  assign new_n_n314_ = ~new_n_n2172_;
  assign new_n_n306_ = ~new_n_n2178_;
  assign new_n_n297_ = ~new_n_n2188_;
  assign new_n_n289_ = ~new_n_n2195_;
  assign new_n_n263_ = ~new_nb4_;
  assign new_n_n255_ = ~new_n_n2230_;
  assign new_n_n246_ = ~new_n_n2235_;
  assign new_n_n222_ = ~new_n_n2258_;
  assign new_n_n214_ = ~new_n_n2265_;
  assign new_n_n205_ = ~new_n_n2276_;
  assign new_n_n196_ = ~new_nina0_;
  assign new_n_n170_ = ~new_nina2_;
  assign new_n_n162_ = ~new_nb3_;
  assign new_n_n1601_ = ~new_ninc13_;
  assign new_n_n121_ = ~new_n_n2360_;
  assign new_n_n113_ = ~new_n_n2363_;
  assign new_n_n104_ = ~new_n_n2159_;
  assign new_n_n2459_ = new_n_n1608_ | new_n_n1715_;
  assign new_n_n1584_ = new_n_n28_ & new_n_n1714_;
  assign new_n_n2442_ = new_n_n1581_ | new_n_n35_;
  assign new_n_n1562_ = new_n_n90_ & new_n_n80_;
  assign new_n_n2381_ = new_n_n1555_ | new_n_n1557_ | new_n_n1556_ | new_n_n1358_;
  assign new_n_n1552_ = new_n_n93_ & new_n_n94_;
  assign new_n_n1528_ = new_n_n129_ & new_n_n1715_;
  assign new_n_n2341_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n135_;
  assign new_n_n2336_ = new_n_n1516_ | new_n_n1518_ | new_n_n1517_ | new_n_n1358_;
  assign new_n_n1501_ = new_n_n104_ & new_n_n162_;
  assign new_n_n2310_ = new_n_n1495_ | new_n_n819_;
  assign new_n_n2299_ = new_n_n1715_ | new_n_n820_ | new_n_n781_;
  assign new_n_n1478_ = new_n_n183_ & new_n_n1714_;
  assign new_n_n2289_ = new_n_n189_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n1454_ = new_n_n1699_ & new_n_n728_;
  assign new_n_n2263_ = new_n_n1448_ | new_n_n819_;
  assign new_n_n2257_ = new_n_n1443_ | new_n_n1444_;
  assign new_n_n1439_ = new_n_n1714_ & new_n_n226_;
  assign new_n_n1437_ = new_n_n228_ & new_n_n229_;
  assign new_n_n1433_ = new_n_n2159_ & new_nb6_;
  assign new_n_n2242_ = new_n_n238_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2221_ = new_n_n260_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2217_ = new_n_n1688_ & new_n_n695_;
  assign new_n_n1397_ = new_n_n271_ & new_n_n272_;
  assign new_n_n1392_ = new_n_n1714_ & new_n_n276_;
  assign new_n_n1380_ = new_n_n1714_ & new_n_n290_;
  assign new_n_n2163_ = new_n_n1349_ | new_n_n1351_ | new_n_n1350_ | new_n_n893_;
  assign new_n_n2000_ = new_n_n1168_ | new_n_n1170_ | new_n_n1169_ | new_n_n893_;
  assign new_n_n1165_ = new_n_n831_ & new_n_n627_;
  assign new_n_n1117_ = new_n_n572_ & new_n_n571_;
  assign new_n_n1954_ = new_n_n1109_ | new_n_n1111_ | new_n_n1110_ | new_n_n893_;
  assign new_n_n1067_ = new_n_n833_ & new_n_n628_;
  assign new_n_n1061_ = new_n_n635_ & new_n_n1676_;
  assign new_n_n1882_ = new_n_n1035_ | new_n_n668_;
  assign new_n_n1877_ = new_n_n2226_ | new_n_n1687_;
  assign new_n_n1024_ = new_n_n676_ & new_n_n640_;
  assign new_n_n1002_ = new_n_n699_ & new_n_n702_;
  assign new_n_n1854_ = new_n_n1724_ | new_n_n703_;
  assign new_n_n1843_ = new_n_n1071_ | new_n_n957_;
  assign new_n_n1837_ = new_n_n973_ | new_n_n913_ | new_n_n974_ | new_n_n975_;
  assign new_n_n969_ = new_n_n728_ & new_n_n729_;
  assign new_n_n967_ = new_n_n742_ & new_n_n741_;
  assign new_n_n1812_ = new_n_n920_ | new_n_n879_ | new_n_n951_ | new_n_n952_;
  assign new_n_n947_ = new_n_n853_ & new_n_n1704_;
  assign new_n_n941_ = new_n_n734_ & new_n_n772_;
  assign new_n_n935_ = new_n_n774_ & new_n_n737_;
  assign new_n_n933_ = new_n_n773_ & new_n_n774_;
  assign new_n_n927_ = new_n_n781_ & new_n_n782_;
  assign new_n_n922_ = new_n_n833_ & new_n_n787_;
  assign new_n_n1782_ = new_n_n794_ | new_n_n795_;
  assign new_n_n901_ = new_n_n848_ & new_n_n1729_;
  assign new_n_n1765_ = new_n_n894_ | new_n_n895_;
  assign new_n_n1760_ = new_n_n889_ | new_n_n821_;
  assign new_n_n883_ = new_n_n790_ & new_n_n1720_;
  assign new_n_n1746_ = new_n_n866_ | new_n_n867_;
  assign new_no0_ = new_n_n861_ | new_n_n854_;
  assign new_n_n1731_ = ~new_n_n2479_;
  assign new_n_n849_ = ~new_n_n1728_;
  assign new_n_n846_ = ~new_n_n1745_;
  assign new_n_n1722_ = ~new_n_n2392_;
  assign new_n_n832_ = ~new_n_n1686_;
  assign new_n_n823_ = ~new_n_n1759_;
  assign new_n_n782_ = ~new_n_n1794_;
  assign new_n_n771_ = ~new_n_n1706_;
  assign new_n_n1705_ = ~new_n_n2304_;
  assign new_n_n761_ = ~new_n_n1814_;
  assign new_n_n752_ = ~new_n_n1821_;
  assign new_n_n741_ = ~new_n_n1825_;
  assign new_n_n699_ = ~new_n_n1858_;
  assign new_n_n692_ = ~new_n_n1845_;
  assign new_n_n690_ = ~new_n_n1636_;
  assign new_n_n680_ = ~new_n_n1872_;
  assign new_n_n671_ = ~new_n_n1882_;
  assign new_n_n662_ = ~new_n_n1890_;
  assign new_n_n618_ = ~new_n_n1925_;
  assign new_n_n608_ = ~new_n_n1738_;
  assign new_n_n1668_ = ~new_n_n1945_;
  assign new_n_n588_ = ~new_n_n1918_;
  assign new_n_n579_ = ~new_n_n1665_;
  assign new_n_n537_ = ~new_n_n1990_;
  assign new_n_n528_ = ~new_n_n2001_;
  assign new_n_n504_ = ~new_n_n2017_;
  assign new_n_n1650_ = ~new_n_n2029_;
  assign new_n_n448_ = ~new_n_n2068_;
  assign new_n_n438_ = ~new_n_n2074_;
  assign new_n_n412_ = ~new_n_n1632_;
  assign new_n_n396_ = ~new_n_n2104_;
  assign new_n_n369_ = ~new_n_n2125_;
  assign new_n_n360_ = ~new_n_n2137_;
  assign new_n_n313_ = ~new_nb9_;
  assign new_n_n303_ = ~new_n_n2181_;
  assign new_n_n282_ = ~new_nina11_;
  assign new_n_n273_ = ~new_n_n2211_;
  assign new_n_n221_ = ~new_n_n2259_;
  assign new_n_n211_ = ~new_n_n2045_;
  assign new_n_n200_ = ~new_n_n2283_;
  assign new_n_n190_ = ~new_n_n2288_;
  assign new_n_n180_ = ~new_n_n2301_;
  assign new_n_n129_ = ~new_nina13_;
  assign new_n_n118_ = ~new_n_n2359_;
  assign new_n_n108_ = ~new_n_n2376_;
  assign new_n_n97_ = ~new_nina15_;
  assign new_n_n8_ = ~new_n_n2477_;
  assign new_n_n1587_ = new_n_n21_ & new_n_n840_;
  assign new_n_n2450_ = new_n_n29_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2443_ = new_n_n840_ | new_n_n36_;
  assign new_n_n1557_ = new_n_n815_ & new_n_n1599_;
  assign new_n_n2376_ = new_n_n1552_ | new_n_n819_;
  assign new_n_n1527_ = new_n_n129_ & new_n_n1601_;
  assign new_n_n2342_ = new_n_n1602_ | new_n_n1716_;
  assign new_n_n2315_ = new_n_n1498_ | new_n_n1500_ | new_n_n1499_ | new_n_n1358_;
  assign new_n_n1496_ = new_n_n1714_ & new_n_n165_;
  assign new_n_n2298_ = new_n_n1481_ | new_n_n1482_;
  assign new_n_n1479_ = new_n_n79_ & new_n_n184_;
  assign new_n_n2288_ = new_n_n815_ | new_n_n1713_ | new_n_n1717_;
  assign new_n_n2268_ = new_n_n1451_ | new_n_n1453_ | new_n_n1452_ | new_n_n1358_;
  assign new_n_n1449_ = new_n_n1714_ & new_n_n214_;
  assign new_n_n1444_ = new_n_n2159_ & new_nb7_;
  assign new_n_n2252_ = new_n_n1438_ | new_n_n1439_;
  assign new_n_n2250_ = new_n_n1608_ | new_n_n1716_;
  assign new_n_n2245_ = new_n_n1432_ | new_n_n1433_;
  assign new_n_n2241_ = new_n_n815_ | new_n_n1713_ | new_n_n1680_;
  assign new_nb4_ = new_n_n261_ & new_n_n262_;
  assign new_n_n2218_ = new_n_n265_ | new_n_n264_;
  assign new_n_n2210_ = new_n_n1396_ | new_n_n273_;
  assign new_n_n2205_ = new_n_n1391_ | new_n_n1392_;
  assign new_n_n2192_ = new_n_n1379_ | new_n_n819_;
  assign new_n_n2170_ = new_n_n815_ | new_n_n1713_ | new_n_n1659_;
  assign new_n_n1170_ = new_n_n79_ & new_n_n528_;
  assign new_n_n1995_ = new_n_n1165_ | new_n_n1107_;
  assign new_n_n1116_ = new_n_n572_ & new_n_n1724_;
  assign new_n_n1955_ = new_n_n579_ & new_n_n815_;
  assign new_n_n1066_ = new_n_n629_ & new_n_n628_;
  assign new_n_n1062_ = new_n_n853_ & new_n_n1676_;
  assign new_n_n1035_ = new_n_n669_ & new_n_n670_;
  assign new_n_n1030_ = new_n_n673_ & new_n_n674_;
  assign new_n_n1019_ = new_n_n79_ & new_n_n685_;
  assign new_n_n1001_ = new_n_n699_ & new_n_n434_;
  assign new_n_n994_ = new_n_n703_ & new_n_n1724_;
  assign new_n_n1842_ = new_n_n953_ | new_n_n879_ | new_n_n979_ | new_n_n980_;
  assign new_n_n976_ = new_n_n722_ & new_n_n723_;
  assign new_n_n1832_ = new_n_n770_ | new_n_n1706_;
  assign new_n_n968_ = new_n_n742_ & new_n_n740_;
  assign new_n_n952_ = new_n_n833_ & new_n_n759_;
  assign new_n_n1807_ = new_n_n945_ | new_n_n913_ | new_n_n946_ | new_n_n947_;
  assign new_n_n1801_ = new_n_n940_ | new_n_n735_;
  assign new_n_n936_ = new_n_n774_ & new_n_n1700_;
  assign new_n_n1796_ = new_n_n931_ | new_n_n932_;
  assign new_n_n928_ = new_n_n781_ & new_n_n1714_;
  assign new_n_n921_ = new_n_n760_ & new_n_n787_;
  assign new_n_n1783_ = new_n_n840_ | new_n_n1722_;
  assign new_n_n900_ = new_n_n1728_ & new_n_n849_;
  assign new_n_n1766_ = new_n_n814_ & new_n_n815_;
  assign new_n_n889_ = new_n_n83_ & new_n_n822_;
  assign new_n_n884_ = new_n_n790_ & new_n_n827_;
  assign new_n_n867_ = new_n_n845_ & new_n_n858_;
  assign new_n_n1743_ = new_n_n852_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n856_ = ~new_n_n2391_;
  assign new_n_n1728_ = ~new_nopsel0_;
  assign new_n_n1727_ = ~new_n_n2328_;
  assign new_n_n1723_ = ~new_n_n1750_;
  assign new_n_n831_ = ~new_n_n1719_;
  assign new_n_n824_ = ~new_n_n1695_;
  assign new_n_n781_ = ~new_ninb1_;
  assign new_n_n772_ = ~new_n_n1830_;
  assign new_n_n1704_ = ~new_n_n1811_;
  assign new_n_n762_ = ~new_n_n1812_;
  assign new_n_n751_ = ~new_ninb2_;
  assign new_n_n742_ = ~new_n_n1833_;
  assign new_n_n698_ = ~new_n_n1689_;
  assign new_n_n693_ = ~new_n_n1863_;
  assign new_n_n689_ = ~new_n_n1865_;
  assign new_n_n681_ = ~new_n_n1871_;
  assign new_n_n1682_ = ~new_n_n1881_;
  assign new_n_n663_ = ~new_n_n1630_;
  assign new_n_n617_ = ~new_n_n1926_;
  assign new_n_n609_ = ~new_n_n1932_;
  assign new_n_n604_ = ~new_n_n1672_;
  assign new_n_n587_ = ~new_n_n1947_;
  assign new_n_n580_ = ~new_ninb7_;
  assign new_n_n536_ = ~new_n_n1989_;
  assign new_n_n1653_ = ~new_nind9_;
  assign new_n_n503_ = ~new_n_n2018_;
  assign new_n_n495_ = ~new_n_n2025_;
  assign new_n_n447_ = ~new_n_n2067_;
  assign new_n_n439_ = ~new_n_n2072_;
  assign new_n_n421_ = ~new_n_n2085_;
  assign new_n_n388_ = ~new_n_n2113_;
  assign new_n_n368_ = ~new_n_n2126_;
  assign new_n_n1623_ = ~new_n_n2135_;
  assign new_n_n312_ = ~new_n_n2177_;
  assign new_n_n304_ = ~new_n_n2180_;
  assign new_n_n281_ = ~new_n_n1612_;
  assign new_n_n1611_ = ~new_n_n2210_;
  assign new_n_n220_ = ~new_n_n2260_;
  assign new_n_n212_ = ~new_n_n2268_;
  assign new_n_n191_ = ~new_n_n2287_;
  assign new_n_n189_ = ~new_n_n2290_;
  assign new_n_n181_ = ~new_n_n2296_;
  assign new_n_n128_ = ~new_nb13_;
  assign new_n_n119_ = ~new_n_n2358_;
  assign new_n_n107_ = ~new_n_n2370_;
  assign new_n_n98_ = ~new_n_n2373_;
  assign new_n_n2457_ = new_n_n1586_ | new_n_n22_;
  assign new_n_n2452_ = new_n_n1714_ | new_n_n815_ | new_n_n245_;
  assign new_n_n2444_ = new_n_n34_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2386_ = new_n_n1561_ | new_n_n82_;
  assign new_n_n1553_ = new_n_n1714_ & new_n_n92_;
  assign new_n_n2347_ = new_n_n130_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n1520_ = new_n_n2159_ & new_nb12_;
  assign new_n_n2305_ = new_n_n172_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n1485_ = new_n_n815_ & new_n_n1605_;
  assign new_n_n1482_ = new_n_n1714_ & new_n_n177_;
  assign new_n_n2292_ = new_n_n185_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n1473_ = new_n_n196_ & new_n_n1715_;
  assign new_n_n1453_ = new_n_n815_ & new_n_n1607_;
  assign new_n_n2262_ = new_n_n1607_ | new_n_n1716_;
  assign new_n_n2258_ = new_n_n221_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2253_ = new_n_n1715_ | new_n_n820_ | new_n_n621_;
  assign new_n_n2249_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n230_;
  assign new_n_n2244_ = new_n_n1428_ | new_n_n1430_ | new_n_n1429_ | new_n_n1431_;
  assign new_n_n1426_ = new_n_n245_ & new_n_n1715_;
  assign new_n_n2220_ = new_n_n1406_ | new_n_n1407_;
  assign new_n_n2215_ = new_n_n1400_ | new_n_n1401_;
  assign new_n_n2212_ = new_n_n598_ | new_n_n1670_;
  assign new_n_n2206_ = new_n_n1715_ | new_n_n820_ | new_n_n445_;
  assign new_n_n2202_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n280_;
  assign new_n_n2197_ = new_n_n1382_ | new_n_n1384_ | new_n_n1383_ | new_n_n1358_;
  assign new_nb9_ = new_n_n311_ & new_n_n312_;
  assign new_n_n2050_ = new_n_n1724_ | new_n_n461_;
  assign new_n_n2043_ = new_n_n1211_ | new_n_n468_;
  assign new_n_n1171_ = new_n_n525_ & new_n_n1730_;
  assign new_n_n1166_ = new_n_n690_ & new_n_n1719_;
  assign new_n_n1959_ = new_n_n1116_ | new_n_n913_ | new_n_n1117_ | new_n_n1118_;
  assign new_n_n1112_ = new_n_n578_ & new_n_n1730_;
  assign new_n_n1910_ = new_n_n1060_ | new_n_n913_ | new_n_n1061_ | new_n_n1062_;
  assign new_n_n1881_ = new_n_n1032_ | new_n_n913_ | new_n_n1033_ | new_n_n1034_;
  assign new_n_n1025_ = new_n_n677_ & new_n_n645_;
  assign new_n_n1869_ = new_n_n1017_ | new_n_n1019_ | new_n_n1018_ | new_n_n893_;
  assign new_n_n1850_ = new_n_n987_ | new_n_n989_ | new_n_n988_ | new_n_n893_;
  assign new_n_n984_ = new_n_n831_ & new_n_n829_;
  assign new_n_n980_ = new_n_n833_ & new_n_n717_;
  assign new_n_n974_ = new_n_n724_ & new_n_n1697_;
  assign new_n_n1833_ = new_n_n969_ | new_n_n970_;
  assign new_n_n1824_ = new_n_n967_ | new_n_n968_;
  assign new_n_n951_ = new_n_n760_ & new_n_n759_;
  assign new_n_n945_ = new_n_n766_ & new_n_n1724_;
  assign new_n_n1802_ = new_n_n941_ | new_n_n942_;
  assign new_n_n1797_ = new_n_n935_ | new_n_n936_;
  assign new_n_n932_ = new_n_n351_ & new_n_n775_;
  assign new_n_n1791_ = new_n_n926_ | new_n_n783_;
  assign new_n_n923_ = new_n_n831_ & new_n_n786_;
  assign new_n_n916_ = new_n_n792_ & new_n_n1721_;
  assign new_n_n899_ = new_n_n1728_ & new_n_n1729_;
  assign new_n_n894_ = new_n_n816_ & new_n_n1715_;
  assign new_n_n1762_ = new_n_n1714_ & new_n_n1715_;
  assign new_n_n885_ = new_n_n833_ & new_n_n827_;
  assign new_n_n1753_ = new_n_n877_ | new_n_n879_ | new_n_n878_ | new_n_n880_;
  assign new_n_n1750_ = new_n_n870_ | new_n_n913_ | new_n_n871_ | new_n_n872_;
  assign new_n_n857_ = ~new_n_n1633_;
  assign new_n_n1729_ = ~new_nopsel1_;
  assign new_n_n1726_ = ~new_n_n2285_;
  assign new_n_n839_ = ~new_n_n1722_;
  assign new_n_n834_ = ~new_n_n1755_;
  assign new_n_n825_ = ~new_n_n1708_;
  assign new_n_n783_ = ~new_n_n1792_;
  assign new_n_n773_ = ~new_n_n1797_;
  assign new_n_n769_ = ~new_n_n1703_;
  assign new_n_n759_ = ~new_n_n1813_;
  assign new_n_n753_ = ~new_n_n1819_;
  assign new_n_n743_ = ~new_n_n1824_;
  assign new_n_n700_ = ~new_n_n1692_;
  assign new_n_n694_ = ~new_n_n1861_;
  assign new_n_n688_ = ~new_n_n1866_;
  assign new_n_n678_ = ~new_n_n1683_;
  assign new_n_n673_ = ~new_n_n1879_;
  assign new_n_n1681_ = ~new_n_n1892_;
  assign new_n_n620_ = ~new_n_n1673_;
  assign new_n_n610_ = ~new_n_n1929_;
  assign new_n_n603_ = ~new_n_n1933_;
  assign new_n_n596_ = ~new_n_n1939_;
  assign new_n_n581_ = ~new_n_n1955_;
  assign new_n_n1655_ = ~new_n_n1987_;
  assign new_n_n529_ = ~new_n_n1999_;
  assign new_n_n523_ = ~new_n_n2003_;
  assign new_n_n512_ = ~new_n_n2012_;
  assign new_n_n450_ = ~new_n_n2061_;
  assign new_n_n440_ = ~new_n_n2071_;
  assign new_n_n429_ = ~new_n_n1637_;
  assign new_n_n378_ = ~new_n_n2123_;
  assign new_n_n1625_ = ~new_n_n2131_;
  assign new_n_n361_ = ~new_n_n2134_;
  assign new_n_n294_ = ~new_n_n1613_;
  assign new_n_n284_ = ~new_n_n2200_;
  assign new_n_n274_ = ~new_n_n2044_;
  assign new_n_n219_ = ~new_nina7_;
  assign new_n_n202_ = ~new_n_n2303_;
  assign new_n_n192_ = ~new_n_n2286_;
  assign new_n_n127_ = ~new_n_n2353_;
  assign new_n_n1600_ = ~new_ninc14_;
  assign new_n_n110_ = ~new_n_n1600_;
  assign new_n_n99_ = ~new_n_n2372_;
  assign new_n_n2458_ = new_n_n1714_ | new_n_n815_ | new_n_n232_;
  assign new_n_n2451_ = new_n_n1584_ | new_n_n27_;
  assign new_n_n1582_ = new_n_n33_ & new_n_n1714_;
  assign new_n_n2387_ = new_n_n1716_ | new_n_n820_ | new_n_n1598_ | new_n_n81_;
  assign new_n_n1558_ = new_n_n87_ & new_n_n88_;
  assign new_n_n2340_ = new_n_n136_ & new_n_n815_;
  assign new_n_n1519_ = new_n_n104_ & new_n_n141_;
  assign new_nb2_ = new_n_n173_ & new_n_n174_;
  assign new_n_n2302_ = new_n_n1483_ | new_n_n1485_ | new_n_n1484_ | new_n_n1358_;
  assign new_n_n1481_ = new_n_n1714_ & new_n_n178_;
  assign new_n_n1477_ = new_n_n183_ & new_n_n184_;
  assign new_n_n1472_ = new_n_n196_ & new_n_n1606_;
  assign new_n_n1452_ = new_n_n219_ & new_n_n1715_;
  assign new_n_n1448_ = new_n_n215_ & new_n_n216_;
  assign new_nb7_ = new_n_n222_ & new_n_n223_;
  assign new_n_n2254_ = new_n_n815_ | new_n_n1713_ | new_n_n1673_;
  assign new_n_n2248_ = new_n_n231_ & new_n_n815_;
  assign new_n_n1432_ = new_n_n104_ & new_n_n237_;
  assign new_n_n1425_ = new_n_n245_ & new_n_n1609_;
  assign new_n_n1407_ = new_n_n2159_ & new_nb4_;
  assign new_n_n2216_ = new_n_n1684_ & new_n_n675_;
  assign new_n_n2211_ = new_n_n1397_ | new_n_n270_;
  assign new_n_n2207_ = new_n_n815_ | new_n_n1713_ | new_n_n1644_;
  assign new_n_n2201_ = new_n_n281_ & new_n_n815_;
  assign new_n_n1385_ = new_n_n104_ & new_n_n287_;
  assign new_n_n2179_ = new_n_n1364_ | new_n_n819_;
  assign new_n_n2049_ = new_n_n462_ & new_n_n351_;
  assign new_n_n2044_ = new_n_n1671_ & new_n_n211_;
  assign new_n_n2001_ = new_n_n526_ & new_n_n815_;
  assign new_n_n1996_ = new_n_n1166_ | new_n_n531_;
  assign new_n_n1118_ = new_n_n853_ & new_n_n571_;
  assign new_n_n1113_ = new_n_n576_ & new_n_n577_;
  assign new_n_n1915_ = new_n_n1040_ | new_n_n879_ | new_n_n1066_ | new_n_n1067_;
  assign new_n_n1876_ = new_n_n1029_ | new_n_n644_;
  assign new_ne5_ = new_n_n1023_ | new_n_n1024_;
  assign new_n_n1870_ = new_n_n683_ & new_n_n815_;
  assign new_n_n989_ = new_n_n79_ & new_n_n711_;
  assign new_n_n1845_ = new_n_n984_ | new_n_n925_;
  assign new_n_n979_ = new_n_n718_ & new_n_n717_;
  assign new_n_n975_ = new_n_n853_ & new_n_n1697_;
  assign new_n_n970_ = new_n_n1698_ & new_n_n1699_;
  assign new_n_n1825_ = new_n_n739_ | new_n_n738_;
  assign new_n_n1811_ = new_n_n949_ | new_n_n950_;
  assign new_n_n946_ = new_n_n766_ & new_n_n1704_;
  assign new_n_n942_ = new_n_n734_ & new_n_n1727_;
  assign new_n_n1798_ = new_n_n736_ | new_n_n735_;
  assign new_n_n931_ = new_n_n385_ & new_n_n776_;
  assign new_n_n1792_ = new_n_n1707_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1787_ = new_n_n920_ | new_n_n879_ | new_n_n921_ | new_n_n922_;
  assign new_n_n917_ = new_n_n836_ & new_n_n791_;
  assign new_n_n1769_ = new_n_n897_ | new_n_n898_;
  assign new_n_n895_ = new_n_n815_ & new_n_n1714_;
  assign new_n_n1761_ = new_n_n1717_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1756_ = new_n_n883_ | new_n_n879_ | new_n_n884_ | new_n_n885_;
  assign new_n_n880_ = new_n_n833_ & new_n_n834_;
  assign new_n_n873_ = new_n_n1722_ & new_n_n1731_;
  assign new_n_n1732_ = ~new_n_n2349_;
  assign new_n_n850_ = ~new_n_n1725_;
  assign new_n_n845_ = ~new_n_n1733_;
  assign new_n_n840_ = ~new_n_n1731_;
  assign new_n_n833_ = ~new_n_n1720_;
  assign new_n_n826_ = ~new_n_n1681_;
  assign new_n_n1707_ = ~new_nind1_;
  assign new_n_n774_ = ~new_n_n1800_;
  assign new_n_n768_ = ~new_n_n1805_;
  assign new_n_n760_ = ~new_n_n1788_;
  assign new_n_n1701_ = ~new_nind2_;
  assign new_n_n744_ = ~new_n_n1827_;
  assign new_n_n1691_ = ~new_n_n1742_;
  assign new_n_n695_ = ~new_n_n1687_;
  assign new_n_n687_ = ~new_n_n1869_;
  assign new_n_n679_ = ~new_ne5_;
  assign new_n_n672_ = ~new_n_n1880_;
  assign new_n_n664_ = ~new_n_n1887_;
  assign new_n_n619_ = ~new_n_n1938_;
  assign new_n_n1672_ = ~new_n_n1936_;
  assign new_n_n602_ = ~new_n_n1934_;
  assign new_n_n597_ = ~new_n_n1667_;
  assign new_n_n589_ = ~new_n_n1948_;
  assign new_n_n538_ = ~new_n_n2423_;
  assign new_n_n530_ = ~new_n_n2000_;
  assign new_n_n522_ = ~new_ne10_;
  assign new_n_n513_ = ~new_n_n1982_;
  assign new_n_n449_ = ~new_n_n2065_;
  assign new_n_n441_ = ~new_n_n1643_;
  assign new_n_n1641_ = ~new_npgx3_;
  assign new_n_n371_ = ~new_n_n1628_;
  assign new_n_n370_ = ~new_n_n1624_;
  assign new_n_n362_ = ~new_n_n2132_;
  assign new_n_n1613_ = ~new_ninc10_;
  assign new_n_n285_ = ~new_n_n2199_;
  assign new_n_n283_ = ~new_n_n2201_;
  assign new_n_n210_ = ~new_n_n2270_;
  assign new_n_n201_ = ~new_nb0_;
  assign new_n_n193_ = ~new_n_n2289_;
  assign new_n_n126_ = ~new_n_n2350_;
  assign new_n_n117_ = ~new_n_n2361_;
  assign new_n_n109_ = ~new_n_n2367_;
  assign new_n_n100_ = ~new_n_n2371_;
  assign new_n_n2484_ = new_n_n1596_ | new_n_n0_;
  assign new_n_n2477_ = new_n_n1601_ | new_n_n1715_;
  assign new_n_n2437_ = new_n_n39_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n1577_ = new_n_n46_ & new_n_n840_;
  assign new_n_n2420_ = new_n_n1574_ | new_n_n52_;
  assign new_n_n2412_ = new_n_n59_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n1569_ = new_n_n66_ & new_n_n840_;
  assign new_n_n2395_ = new_n_n1566_ | new_n_n72_;
  assign new_n_n1564_ = new_n_n79_ & new_n_n80_;
  assign new_n_n2365_ = new_n_n110_ & new_n_n815_;
  assign new_n_n1540_ = new_n_n815_ & new_n_n1600_;
  assign new_n_n2355_ = new_n_n2356_ | new_n_n1626_;
  assign new_n_n1531_ = new_n_n2159_ & new_nb13_;
  assign new_n_n1525_ = new_n_n1714_ & new_n_n132_;
  assign new_nb12_ = new_n_n139_ & new_n_n140_;
  assign new_n_n2331_ = new_n_n1513_ | new_n_n819_;
  assign new_n_n1484_ = new_n_n183_ & new_n_n1715_;
  assign new_n_n2295_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n181_;
  assign new_n_n2290_ = new_n_n1472_ | new_n_n1474_ | new_n_n1473_ | new_n_n1358_;
  assign new_n_n2282_ = new_n_n195_ & new_n_n815_;
  assign new_n_n1463_ = new_n_n1726_ & new_n_n1712_;
  assign new_n_n1457_ = new_n_n206_ & new_n_n1706_;
  assign new_n_n2235_ = new_n_n244_ & new_n_n815_;
  assign new_n_n1416_ = new_n_n815_ & new_n_n1610_;
  assign new_n_n2225_ = new_n_n1610_ | new_n_n1716_;
  assign new_n_n2184_ = new_n_n1367_ | new_n_n1369_ | new_n_n1368_ | new_n_n1358_;
  assign new_n_n2038_ = new_n_n1206_ | new_n_n1207_;
  assign new_n_n1201_ = new_n_n480_ & new_n_n481_;
  assign new_n_n1992_ = new_n_n1134_ | new_n_n879_ | new_n_n1159_ | new_n_n1160_;
  assign new_n_n1155_ = new_n_n853_ & new_n_n1656_;
  assign new_n_n1982_ = new_n_n2167_ | new_n_n1617_;
  assign new_n_n1978_ = new_n_n548_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n1973_ = new_n_n1719_ | new_n_n1660_;
  assign new_n_n1951_ = new_n_n1719_ | new_n_n1666_;
  assign new_n_n1102_ = new_n_n833_ & new_n_n587_;
  assign new_n_n1096_ = new_n_n594_ & new_n_n1668_;
  assign new_n_n1935_ = new_n_n2045_ | new_n_n600_;
  assign new_n_n1085_ = new_n_n605_ & new_n_n644_;
  assign new_n_n1079_ = new_n_n351_ & new_n_n615_;
  assign new_n_n1921_ = new_n_n1073_ | new_n_n623_;
  assign new_n_n1916_ = new_n_n1165_ | new_n_n1044_;
  assign new_n_n1055_ = new_n_n650_ & new_n_n606_;
  assign new_n_n1895_ = new_n_n656_ & new_n_n815_;
  assign new_n_n1889_ = new_n_n1043_ | new_n_n985_;
  assign new_n_n1037_ = new_n_n836_ & new_n_n666_;
  assign new_n_n1879_ = new_n_n672_ & new_n_n351_;
  assign new_n_n1873_ = new_n_n1025_ | new_n_n1026_;
  assign new_n_n1020_ = new_n_n682_ & new_n_n1730_;
  assign new_n_n1844_ = new_n_n981_ | new_n_n879_ | new_n_n982_ | new_n_n983_;
  assign new_n_n1840_ = new_n_n840_ | new_n_n795_ | new_n_n1722_ | new_n_n765_;
  assign new_n_n972_ = new_n_n726_ & new_n_n351_;
  assign new_n_n1826_ = new_n_n737_ | new_n_n1700_;
  assign new_n_n1821_ = new_n_n750_ & new_n_n815_;
  assign new_n_n1815_ = new_n_n956_ | new_n_n888_;
  assign new_n_n1784_ = new_n_n916_ | new_n_n917_;
  assign new_n_n1777_ = new_n_n909_ | new_n_n910_;
  assign new_n_n906_ = new_n_n808_ & new_n_n772_;
  assign new_n_n1714_ = ~new_nmusel1_;
  assign new_n_n810_ = ~new_ne1_;
  assign new_n_n1711_ = ~new_n_n2291_;
  assign new_n_n792_ = ~new_n_n1785_;
  assign new_n_n735_ = ~new_n_n1829_;
  assign new_n_n727_ = ~new_n_n1696_;
  assign new_n_n717_ = ~new_n_n1843_;
  assign new_n_n708_ = ~new_n_n1852_;
  assign new_n_n656_ = ~new_n_n1680_;
  assign new_n_n645_ = ~new_n_n1874_;
  assign new_n_n638_ = ~new_n_n1675_;
  assign new_n_n628_ = ~new_n_n1916_;
  assign new_n_n614_ = ~new_n_n1931_;
  assign new_n_n1661_ = ~new_n_n1965_;
  assign new_n_n555_ = ~new_n_n1976_;
  assign new_n_n545_ = ~new_n_n1983_;
  assign new_n_n533_ = ~new_n_n1971_;
  assign new_n_n524_ = ~new_n_n2002_;
  assign new_n_n468_ = ~new_n_n1611_;
  assign new_n_n460_ = ~new_n_n2435_;
  assign new_n_n445_ = ~new_ninb11_;
  assign new_n_n436_ = ~new_n_n1641_;
  assign new_n_n430_ = ~new_n_n1638_;
  assign new_n_n377_ = ~new_n_n2090_;
  assign new_n_n366_ = ~new_n_n2478_;
  assign new_n_n357_ = ~new_ninb14_;
  assign new_n_n1621_ = ~new_n_n2355_;
  assign new_n_n336_ = ~new_n_n2156_;
  assign new_n_n279_ = ~new_n_n2208_;
  assign new_n_n269_ = ~new_n_n2215_;
  assign new_n_n258_ = ~new_nina4_;
  assign new_n_n248_ = ~new_n_n2233_;
  assign new_n_n238_ = ~new_n_n2243_;
  assign new_n_n186_ = ~new_n_n2292_;
  assign new_n_n176_ = ~new_n_n2302_;
  assign new_n_n166_ = ~new_n_n2311_;
  assign new_n_n1603_ = ~new_ninc3_;
  assign new_n_n145_ = ~new_n_n2333_;
  assign new_n_n135_ = ~new_n_n2342_;
  assign new_n_n5_ = ~new_n_n2480_;
  assign new_n_n2485_ = new_n_n1714_ | new_n_n815_ | new_n_n116_;
  assign new_n_n2469_ = new_n_n1590_ | new_n_n12_;
  assign new_n_n2436_ = new_n_n840_ | new_n_n41_;
  assign new_n_n2429_ = new_n_n1577_ | new_n_n45_;
  assign new_n_n1574_ = new_n_n53_ & new_n_n1714_;
  assign new_n_n1572_ = new_n_n58_ & new_n_n1714_;
  assign new_n_n2403_ = new_n_n1605_ | new_n_n1715_;
  assign new_n_n2396_ = new_n_n1714_ | new_n_n815_ | new_n_n196_;
  assign new_n_n1563_ = new_n_n90_ & new_n_n1714_;
  assign new_n_n2371_ = new_n_n99_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n1539_ = new_n_n116_ & new_n_n1715_;
  assign new_n_n1535_ = new_n_n120_ & new_n_n121_;
  assign new_n_n1530_ = new_n_n104_ & new_n_n128_;
  assign new_n_n1526_ = new_n_n1714_ & new_n_n131_;
  assign new_n_n2337_ = new_n_n1519_ | new_n_n1520_;
  assign new_n_n1514_ = new_n_n1714_ & new_n_n145_;
  assign new_n_n1483_ = new_n_n183_ & new_n_n1605_;
  assign new_n_n2296_ = new_n_n1605_ | new_n_n1716_;
  assign new_n_n1474_ = new_n_n815_ & new_n_n1606_;
  assign new_n_n2283_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n194_;
  assign new_n_n1462_ = new_n_n1726_ & new_n_n801_;
  assign new_n_n2273_ = new_n_n1456_ | new_n_n1457_;
  assign new_n_n1427_ = new_n_n815_ & new_n_n1609_;
  assign new_n_n2236_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n243_;
  assign new_n_n1415_ = new_n_n258_ & new_n_n1715_;
  assign new_n_n1411_ = new_n_n254_ & new_n_n255_;
  assign new_n_n2187_ = new_n_n297_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n1207_ = new_n_n506_ & new_n_n1616_;
  assign new_n_n1202_ = new_n_n480_ & new_n_n479_;
  assign new_n_n1160_ = new_n_n833_ & new_n_n494_;
  assign new_n_n1987_ = new_n_n1153_ | new_n_n913_ | new_n_n1154_ | new_n_n1155_;
  assign new_n_n1981_ = new_n_n512_ | new_n_n1616_;
  assign new_n_n1143_ = new_n_n385_ & new_n_n547_;
  assign new_n_n1968_ = new_n_n1103_ | new_n_n879_ | new_n_n1131_ | new_n_n1132_;
  assign new_n_n1950_ = new_n_n1107_ | new_n_n584_;
  assign new_n_n1946_ = new_n_n1068_ | new_n_n879_ | new_n_n1101_ | new_n_n1102_;
  assign new_n_n1095_ = new_n_n594_ & new_n_n1724_;
  assign new_n_n1936_ = new_n_n2251_ | new_n_n1677_;
  assign new_n_n1929_ = new_n_n1084_ | new_n_n606_;
  assign new_n_n1926_ = new_n_n1078_ | new_n_n1079_;
  assign new_n_n1073_ = new_n_n83_ & new_n_n624_;
  assign new_n_n1068_ = new_n_n588_ & new_n_n1720_;
  assign new_n_n1905_ = new_n_n2238_ | new_n_n1734_;
  assign new_n_n1894_ = new_n_n1046_ | new_n_n1048_ | new_n_n1047_ | new_n_n893_;
  assign new_n_n1044_ = new_n_n829_ & new_n_n1719_;
  assign new_n_n1036_ = new_n_n667_ & new_n_n1721_;
  assign new_n_n1880_ = new_n_n1724_ | new_n_n671_;
  assign new_n_n1026_ = new_n_n677_ & new_n_n1679_;
  assign new_no5_ = new_n_n1020_ | new_n_n681_;
  assign new_n_n983_ = new_n_n833_ & new_n_n715_;
  assign new_n_n977_ = new_n_n720_ & new_n_n1721_;
  assign new_n_n971_ = new_n_n726_ & new_n_n727_;
  assign new_n_n1827_ = new_n_n733_ | new_n_n738_;
  assign new_n_n1820_ = new_n_n959_ | new_n_n961_ | new_n_n960_ | new_n_n893_;
  assign new_n_n957_ = new_n_n826_ & new_n_n1719_;
  assign new_n_n924_ = new_n_n828_ & new_n_n1719_;
  assign new_n_n910_ = new_n_n798_ & new_n_n351_;
  assign new_n_n1771_ = new_n_n905_ | new_n_n906_;
  assign new_n_n1713_ = ~new_nmusel3_;
  assign new_n_n811_ = ~new_n_n1769_;
  assign new_n_n800_ = ~new_n_n1775_;
  assign new_n_n793_ = ~new_n_n1782_;
  assign new_n_n734_ = ~new_n_n1739_;
  assign new_n_n1697_ = ~new_n_n1841_;
  assign new_n_n1695_ = ~new_n_n1848_;
  assign new_n_n709_ = ~new_n_n1694_;
  assign new_n_n655_ = ~new_n_n1907_;
  assign new_n_n646_ = ~new_n_n1900_;
  assign new_n_n637_ = ~new_n_n1908_;
  assign new_n_n629_ = ~new_n_n1889_;
  assign new_n_n605_ = ~new_n_n1737_;
  assign new_n_n1664_ = ~new_n_n1959_;
  assign new_n_n554_ = ~new_n_n1975_;
  assign new_n_n546_ = ~new_n_n1656_;
  assign new_n_n1654_ = ~new_n_n1998_;
  assign new_n_n525_ = ~new_n_n2016_;
  assign new_n_n1647_ = ~new_n_n2192_;
  assign new_n_n1645_ = ~new_n_n2051_;
  assign new_n_n444_ = ~new_n_n1644_;
  assign new_n_n1642_ = ~new_n_n2466_;
  assign new_n_n1635_ = ~new_n_n2386_;
  assign new_n_n387_ = ~new_n_n2114_;
  assign new_n_n365_ = ~new_n_n2130_;
  assign new_n_n358_ = ~new_n_n2138_;
  assign new_n_n346_ = ~new_n_n2143_;
  assign new_n_n337_ = ~new_ng3_;
  assign new_n_n278_ = ~new_n_n2205_;
  assign new_n_n270_ = ~new_n_n2212_;
  assign new_n_n257_ = ~new_n_n1610_;
  assign new_n_n249_ = ~new_n_n2236_;
  assign new_n_n229_ = ~new_n_n2255_;
  assign new_n_n185_ = ~new_n_n2293_;
  assign new_n_n177_ = ~new_n_n2300_;
  assign new_n_n165_ = ~new_n_n2312_;
  assign new_n_n156_ = ~new_n_n1603_;
  assign new_n_n144_ = ~new_n_n2334_;
  assign new_n_n136_ = ~new_n_n1602_;
  assign new_n_n6_ = ~new_n_n1597_;
  assign new_n_n2486_ = new_n_n1600_ | new_n_n1715_;
  assign new_n_n2462_ = new_n_n19_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2435_ = new_n_n1579_ | new_n_n40_;
  assign new_n_n2427_ = new_n_n1714_ | new_n_n815_ | new_n_n308_;
  assign new_n_n2422_ = new_n_n1615_ | new_n_n1715_;
  assign new_n_n2413_ = new_n_n1572_ | new_n_n57_;
  assign new_n_n2402_ = new_n_n1714_ | new_n_n815_ | new_n_n183_;
  assign new_n_n2394_ = new_n_n74_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2389_ = new_n_n815_ & new_n_n78_;
  assign new_nb15_ = new_n_n100_ & new_n_n101_;
  assign new_n_n1545_ = new_n_n79_ & new_n_n111_;
  assign new_n_n2356_ = new_n_n1535_ | new_n_n819_;
  assign new_n_n2348_ = new_n_n1527_ | new_n_n1529_ | new_n_n1528_ | new_n_n1358_;
  assign new_n_n1524_ = new_n_n133_ & new_n_n134_;
  assign new_n_n1521_ = new_n_n142_ & new_n_n137_;
  assign new_n_n1509_ = new_n_n157_ & new_n_n1603_;
  assign new_n_n2319_ = new_n_n156_ & new_n_n815_;
  assign new_n_n2301_ = new_n_n176_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2293_ = new_n_n1477_ | new_n_n1479_ | new_n_n1478_ | new_n_n893_;
  assign new_n_n1476_ = new_n_n2159_ & new_nb1_;
  assign new_n_n1468_ = new_n_n79_ & new_n_n197_;
  assign new_n_n1464_ = new_n_n104_ & new_n_n201_;
  assign new_n_n1458_ = new_n_n204_ & new_n_n205_;
  assign new_nb6_ = new_n_n235_ & new_n_n236_;
  assign new_n_n1421_ = new_n_n79_ & new_n_n246_;
  assign new_n_n1417_ = new_n_n104_ & new_n_n250_;
  assign new_n_n2226_ = new_n_n1411_ | new_n_n819_;
  assign new_n_n1197_ = new_n_n79_ & new_n_n489_;
  assign new_n_n1191_ = new_n_n494_ & new_n_n493_;
  assign new_n_n1159_ = new_n_n533_ & new_n_n494_;
  assign new_n_n1153_ = new_n_n539_ & new_n_n1724_;
  assign new_n_n1150_ = new_n_n1735_ & new_n_n1658_;
  assign new_n_n1144_ = new_n_n351_ & new_n_n546_;
  assign new_n_n1127_ = new_n_n1661_ & new_n_n565_;
  assign new_n_n1107_ = new_n_n758_ & new_n_n1719_;
  assign new_n_n1945_ = new_n_n1099_ | new_n_n1100_;
  assign new_n_n1941_ = new_n_n1095_ | new_n_n913_ | new_n_n1096_ | new_n_n1097_;
  assign new_n_n1091_ = new_n_n598_ & new_n_n599_;
  assign new_n_n1084_ = new_n_n607_ & new_n_n608_;
  assign new_n_n1925_ = new_n_n617_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n1074_ = new_n_n621_ & new_n_n622_;
  assign new_n_n1069_ = new_n_n588_ & new_n_n626_;
  assign new_n_n1904_ = new_n_n695_ | new_n_n1688_;
  assign new_ne6_ = new_n_n1052_ | new_n_n1053_;
  assign new_n_n1890_ = new_n_n1044_ | new_n_n661_;
  assign new_n_n1884_ = new_n_n1691_ | new_n_n1692_;
  assign new_n_n1031_ = new_n_n673_ & new_n_n351_;
  assign new_n_n1027_ = new_n_n675_ & new_n_n859_;
  assign new_n_n1871_ = new_n_n680_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n1864_ = new_n_n1014_ | new_n_n957_;
  assign new_n_n1008_ = new_n_n836_ & new_n_n693_;
  assign new_n_n982_ = new_n_n692_ & new_n_n715_;
  assign new_n_n1838_ = new_n_n976_ | new_n_n721_;
  assign new_n_n1835_ = new_n_n725_ & new_n_n351_;
  assign new_n_n1828_ = new_n_n732_ | new_n_n740_;
  assign new_no3_ = new_n_n962_ | new_n_n748_;
  assign new_n_n1816_ = new_n_n957_ | new_n_n755_;
  assign new_n_n929_ = new_n_n79_ & new_n_n782_;
  assign new_n_n1779_ = new_n_n1724_ | new_n_n796_;
  assign new_n_n1772_ = new_n_n804_ | new_n_n803_;
  assign new_n_n819_ = ~new_n_n1716_;
  assign new_n_n808_ = ~new_n_n1773_;
  assign new_n_n801_ = ~new_n_n1711_;
  assign new_n_n794_ = ~new_n_n1783_;
  assign new_n_n780_ = ~new_n_n1707_;
  assign new_n_n733_ = ~new_n_n1828_;
  assign new_n_n725_ = ~new_n_n1836_;
  assign new_n_n719_ = ~new_n_n1844_;
  assign new_n_n710_ = ~new_ninb3_;
  assign new_n_n1690_ = ~new_n_n1935_;
  assign new_n_n1686_ = ~new_n_n1867_;
  assign new_n_n654_ = ~new_n_n1896_;
  assign new_n_n644_ = ~new_n_n1904_;
  assign new_n_n639_ = ~new_n_n1679_;
  assign new_n_n630_ = ~new_n_n1917_;
  assign new_n_n616_ = ~new_ne7_;
  assign new_n_n606_ = ~new_n_n1905_;
  assign new_n_n571_ = ~new_n_n1967_;
  assign new_n_n563_ = ~new_n_n1617_;
  assign new_n_n547_ = ~new_ne9_;
  assign new_n_n535_ = ~new_n_n1992_;
  assign new_n_n526_ = ~new_n_n1653_;
  assign new_n_n488_ = ~new_ninb10_;
  assign new_n_n477_ = ~new_n_n2039_;
  assign new_n_n1644_ = ~new_nind11_;
  assign new_n_n437_ = ~new_n_n2078_;
  assign new_n_n413_ = ~new_ne13_;
  assign new_n_n1630_ = ~new_n_n2108_;
  assign new_n_n367_ = ~new_n_n2128_;
  assign new_n_n1622_ = ~new_nind14_;
  assign new_n_n330_ = ~new_n_n2154_;
  assign new_n_n321_ = ~new_nina8_;
  assign new_n_n1612_ = ~new_ninc11_;
  assign new_n_n271_ = ~new_n_n2213_;
  assign new_n_n1610_ = ~new_ninc4_;
  assign new_n_n240_ = ~new_n_n2240_;
  assign new_n_n230_ = ~new_n_n2250_;
  assign new_n_n188_ = ~new_nb1_;
  assign new_n_n178_ = ~new_n_n2299_;
  assign new_n_n164_ = ~new_n_n2313_;
  assign new_n_n154_ = ~new_n_n2326_;
  assign new_n_n147_ = ~new_n_n2335_;
  assign new_n_n137_ = ~new_n_n2340_;
  assign new_n_n1597_ = ~new_n_n2483_;
  assign new_n_n1579_ = new_n_n41_ & new_n_n840_;
  assign new_n_n2428_ = new_n_n1614_ | new_n_n1715_;
  assign new_n_n2421_ = new_n_n1714_ | new_n_n815_ | new_n_n321_;
  assign new_n_n2414_ = new_n_n1714_ | new_n_n815_ | new_n_n157_;
  assign new_n_n2401_ = new_n_n1568_ | new_n_n67_;
  assign new_n_n1566_ = new_n_n73_ & new_n_n1714_;
  assign new_n_n2388_ = new_n_n1562_ | new_n_n1564_ | new_n_n1563_ | new_n_n893_;
  assign new_n_n2370_ = new_n_n1547_ | new_n_n1548_;
  assign new_n_n2364_ = new_n_n1543_ | new_n_n1545_ | new_n_n1544_ | new_n_n893_;
  assign new_n_n2361_ = new_n_n1538_ | new_n_n1540_ | new_n_n1539_ | new_n_n1358_;
  assign new_n_n1529_ = new_n_n815_ & new_n_n1601_;
  assign new_n_n2343_ = new_n_n1524_ | new_n_n819_;
  assign new_n_n2338_ = new_n_n138_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2326_ = new_n_n150_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2320_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n155_;
  assign new_n_n2300_ = new_n_n815_ | new_n_n1713_ | new_n_n1707_;
  assign new_n_n2294_ = new_n_n182_ & new_n_n815_;
  assign new_n_n1475_ = new_n_n104_ & new_n_n188_;
  assign new_n_n2281_ = new_n_n1466_ | new_n_n1468_ | new_n_n1467_ | new_n_n893_;
  assign new_n_n2278_ = new_n_n1460_ | new_n_n1462_ | new_n_n1461_ | new_n_n1463_;
  assign new_n_n1459_ = new_n_n204_ & new_n_n735_;
  assign new_n_n2251_ = new_n_n1437_ | new_n_n819_;
  assign new_n_n2234_ = new_n_n1419_ | new_n_n1421_ | new_n_n1420_ | new_n_n893_;
  assign new_n_n2231_ = new_n_n1414_ | new_n_n1416_ | new_n_n1415_ | new_n_n1358_;
  assign new_n_n1412_ = new_n_n1714_ & new_n_n253_;
  assign new_n_n1196_ = new_n_n488_ & new_n_n1714_;
  assign new_n_n1192_ = new_n_n833_ & new_n_n493_;
  assign new_n_n1991_ = new_n_n1157_ | new_n_n1158_;
  assign new_n_n1154_ = new_n_n539_ & new_n_n1656_;
  assign new_n_n1149_ = new_n_n543_ & new_n_n860_;
  assign new_n_n1979_ = new_n_n1143_ | new_n_n1144_;
  assign new_n_n1960_ = new_n_n1119_ | new_n_n1120_;
  assign new_n_n1949_ = new_n_n1106_ | new_n_n1044_;
  assign new_n_n1101_ = new_n_n588_ & new_n_n587_;
  assign new_n_n1097_ = new_n_n853_ & new_n_n1668_;
  assign new_n_n1092_ = new_n_n1669_ & new_n_n1670_;
  assign new_n_n1928_ = new_n_n610_ | new_n_n609_;
  assign new_n_n1078_ = new_n_n385_ & new_n_n616_;
  assign new_n_n1922_ = new_n_n1673_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1070_ = new_n_n833_ & new_n_n626_;
  assign new_n_n1903_ = new_n_n640_ | new_n_n606_;
  assign new_n_n1054_ = new_n_n650_ & new_n_n647_;
  assign new_n_n1049_ = new_n_n655_ & new_n_n1730_;
  assign new_n_n1883_ = new_n_n669_ | new_n_n670_;
  assign new_n_n1878_ = new_n_n1030_ | new_n_n1031_;
  assign new_n_n1874_ = new_n_n644_ | new_n_n1690_;
  assign new_n_n1021_ = new_n_n385_ & new_n_n679_;
  assign new_n_n1014_ = new_n_n831_ & new_n_n788_;
  assign new_n_n1860_ = new_n_n1007_ | new_n_n1008_;
  assign new_n_n981_ = new_n_n692_ & new_n_n1720_;
  assign new_n_n1839_ = new_n_n722_ | new_n_n723_;
  assign new_n_n1834_ = new_n_n971_ | new_n_n972_;
  assign new_n_n1829_ = new_n_n801_ | new_n_n1712_;
  assign new_n_n962_ = new_n_n749_ & new_n_n1730_;
  assign new_n_n1817_ = new_n_n1719_ | new_n_n1702_;
  assign new_n_n934_ = new_n_n773_ & new_n_n732_;
  assign new_n_n1778_ = new_n_n797_ & new_n_n351_;
  assign new_n_n907_ = new_n_n801_ & new_n_n802_;
  assign new_n_n818_ = ~new_n_n1766_;
  assign new_n_n809_ = ~new_n_n1710_;
  assign new_n_n1712_ = ~new_n_n2297_;
  assign new_n_n795_ = ~new_n_n2398_;
  assign new_n_n770_ = ~new_n_n1705_;
  assign new_n_n732_ = ~new_n_n1801_;
  assign new_n_n726_ = ~new_n_n1835_;
  assign new_n_n718_ = ~new_n_n1815_;
  assign new_n_n711_ = ~new_n_n1851_;
  assign new_n_n697_ = ~new_n_n1690_;
  assign new_n_n691_ = ~new_n_n1862_;
  assign new_n_n653_ = ~new_n_n1897_;
  assign new_n_n1679_ = ~new_n_n1877_;
  assign new_n_n1676_ = ~new_n_n1914_;
  assign new_n_n631_ = ~new_n_n1915_;
  assign new_n_n615_ = ~new_n_n1668_;
  assign new_n_n607_ = ~new_n_n1930_;
  assign new_n_n1663_ = ~new_n_n2417_;
  assign new_n_n564_ = ~new_n_n1657_;
  assign new_n_n556_ = ~new_n_n1973_;
  assign new_n_n534_ = ~new_n_n1994_;
  assign new_n_n527_ = ~new_ninb9_;
  assign new_n_n487_ = ~new_n_n1648_;
  assign new_n_n478_ = ~new_n_n2036_;
  assign new_n_n446_ = ~new_n_n2069_;
  assign new_n_n1643_ = ~new_n_n2073_;
  assign new_n_n405_ = ~new_n_n2098_;
  assign new_n_n1631_ = ~new_n_n2097_;
  assign new_n_n1624_ = ~new_n_n2127_;
  assign new_n_n359_ = ~new_n_n2136_;
  assign new_n_n1617_ = ~new_n_n2158_;
  assign new_n_n322_ = ~new_n_n2164_;
  assign new_n_n280_ = ~new_n_n2203_;
  assign new_n_n272_ = ~new_n_n2214_;
  assign new_n_n247_ = ~new_n_n2234_;
  assign new_n_n239_ = ~new_n_n2241_;
  assign new_n_n1608_ = ~new_ninc6_;
  assign new_n_n187_ = ~new_n_n2295_;
  assign new_n_n179_ = ~new_n_n2298_;
  assign new_n_n163_ = ~new_n_n2315_;
  assign new_n_n155_ = ~new_n_n2321_;
  assign new_n_n146_ = ~new_n_n2332_;
  assign new_n_n138_ = ~new_n_n2339_;
  assign new_n_n7_ = ~new_n_n2476_;
  assign new_n_n2479_ = new_n_n5_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n1591_ = new_n_n11_ & new_n_n840_;
  assign new_n_n2463_ = new_n_n1588_ | new_n_n17_;
  assign new_n_n2434_ = new_n_n1613_ | new_n_n1715_;
  assign new_n_n1576_ = new_n_n48_ & new_n_n1714_;
  assign new_n_n2417_ = new_n_n1573_ | new_n_n55_;
  assign new_n_n2409_ = new_n_n1604_ | new_n_n1715_;
  assign new_n_n1570_ = new_n_n63_ & new_n_n1714_;
  assign new_n_n2398_ = new_n_n1567_ | new_n_n70_;
  assign new_npgx3_ = new_n_n77_ & new_n_n1731_ & new_n_n856_ & new_n_n456_;
  assign new_n_n2382_ = new_n_n1558_ | new_n_n1559_;
  assign new_n_n1554_ = new_n_n1714_ & new_n_n91_;
  assign new_n_n1548_ = new_n_n2159_ & new_nb15_;
  assign new_n_n1543_ = new_n_n116_ & new_n_n111_;
  assign new_n_n2359_ = new_n_n815_ | new_n_n1713_ | new_n_n1622_;
  assign new_n_n2351_ = new_n_n1532_ | new_n_n1534_ | new_n_n1533_ | new_n_n893_;
  assign new_n_n2346_ = new_n_n815_ | new_n_n1713_ | new_n_n1629_;
  assign new_n_n1523_ = new_n_n79_ & new_n_n137_;
  assign new_n_n2333_ = new_n_n1715_ | new_n_n820_ | new_n_n418_;
  assign new_n_n1511_ = new_n_n815_ & new_n_n1603_;
  assign new_n_n2321_ = new_n_n1603_ | new_n_n1716_;
  assign new_n_n2318_ = new_n_n1503_ | new_n_n1505_ | new_n_n1504_ | new_n_n893_;
  assign new_n_n1499_ = new_n_n170_ & new_n_n1715_;
  assign new_n_n2308_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n168_;
  assign new_n_n2303_ = new_n_n1486_ | new_n_n1488_ | new_n_n1487_ | new_n_n1489_;
  assign new_n_n2285_ = new_n_n1469_ | new_n_n819_;
  assign new_n_n2279_ = new_n_n1464_ | new_n_n1465_;
  assign new_n_n2274_ = new_n_n1458_ | new_n_n1459_;
  assign new_n_n2256_ = new_n_n1440_ | new_n_n1442_ | new_n_n1441_ | new_n_n1358_;
  assign new_n_n2232_ = new_n_n1417_ | new_n_n1418_;
  assign new_n_n1413_ = new_n_n1714_ & new_n_n252_;
  assign new_n_n2022_ = new_n_n569_ | new_n_n538_ | new_n_n1663_;
  assign new_n_n1181_ = new_n_n504_ & new_n_n351_;
  assign new_n_n1158_ = new_n_n836_ & new_n_n534_;
  assign new_n_n1139_ = new_n_n552_ & new_n_n553_;
  assign new_n_n1134_ = new_n_n533_ & new_n_n1720_;
  assign new_n_n1128_ = new_n_n563_ & new_n_n564_;
  assign new_n_n1961_ = new_n_n1730_ | new_n_n853_;
  assign new_n_n1106_ = new_n_n831_ & new_n_n690_;
  assign new_n_n1099_ = new_n_n590_ & new_n_n1721_;
  assign new_n_n1938_ = new_n_n1093_ | new_n_n1094_;
  assign new_n_n1089_ = new_n_n608_ & new_n_n606_;
  assign new_n_n1931_ = new_n_n1087_ | new_n_n609_;
  assign new_ne7_ = new_n_n1080_ | new_n_n1081_;
  assign new_n_n1076_ = new_n_n79_ & new_n_n622_;
  assign new_n_n1917_ = new_n_n1068_ | new_n_n879_ | new_n_n1069_ | new_n_n1070_;
  assign new_n_n1063_ = new_n_n633_ & new_n_n634_;
  assign new_n_n1902_ = new_n_n641_ | new_n_n266_;
  assign new_n_n1052_ = new_n_n649_ & new_n_n650_;
  assign new_n_n1046_ = new_n_n657_ & new_n_n658_;
  assign new_n_n1041_ = new_n_n629_ & new_n_n662_;
  assign new_n_n1034_ = new_n_n853_ & new_n_n1683_;
  assign new_n_n1875_ = new_n_n1027_ | new_n_n1028_;
  assign new_n_n1022_ = new_n_n351_ & new_n_n678_;
  assign new_n_n1865_ = new_n_n1015_ | new_n_n688_;
  assign new_n_n1009_ = new_n_n692_ & new_n_n691_;
  assign new_n_n1007_ = new_n_n694_ & new_n_n1721_;
  assign new_n_n999_ = new_n_n568_ & new_n_n434_;
  assign new_n_n993_ = new_n_n705_ & new_n_n351_;
  assign new_n_n1848_ = new_n_n986_ | new_n_n712_;
  assign new_n_n963_ = new_n_n385_ & new_n_n746_;
  assign new_n_n958_ = new_n_n83_ & new_n_n754_;
  assign new_n_n1800_ = new_n_n938_ | new_n_n939_;
  assign new_n_n912_ = new_n_n796_ & new_n_n1710_;
  assign new_n_n908_ = new_n_n1711_ & new_n_n1712_;
  assign new_n_n817_ = ~new_ninb0_;
  assign new_n_n806_ = ~new_n_n1774_;
  assign new_n_n798_ = ~new_n_n1778_;
  assign new_n_n1708_ = ~new_n_n1791_;
  assign new_n_n764_ = ~new_n_n1810_;
  assign new_n_n731_ = ~new_n_n1700_;
  assign new_n_n1696_ = ~new_n_n1837_;
  assign new_n_n714_ = ~new_n_n1847_;
  assign new_n_n704_ = ~new_n_n1854_;
  assign new_n_n683_ = ~new_n_n1685_;
  assign new_n_n674_ = ~new_n_n1682_;
  assign new_n_n652_ = ~new_ne6_;
  assign new_n_n642_ = ~new_n_n1677_;
  assign new_n_n1675_ = ~new_n_n1910_;
  assign new_n_n625_ = ~new_n_n1920_;
  assign new_n_n598_ = ~new_n_n1669_;
  assign new_n_n591_ = ~new_n_n1943_;
  assign new_n_n1665_ = ~new_nind7_;
  assign new_n_n1662_ = ~new_n_n2055_;
  assign new_n_n561_ = ~new_n_n1968_;
  assign new_n_n552_ = ~new_ninb8_;
  assign new_n_n1657_ = ~new_n_n2167_;
  assign new_n_n517_ = ~new_n_n2005_;
  assign new_n_n506_ = ~new_n_n2013_;
  assign new_n_n497_ = ~new_n_n2026_;
  assign new_n_n489_ = ~new_n_n2032_;
  assign new_n_n486_ = ~new_n_n2048_;
  assign new_n_n475_ = ~new_n_n2041_;
  assign new_n_n465_ = ~new_n_n2047_;
  assign new_n_n456_ = ~new_n_n2416_;
  assign new_n_n431_ = ~new_n_n1640_;
  assign new_n_n423_ = ~new_n_n2062_;
  assign new_n_n415_ = ~new_n_n2087_;
  assign new_n_n406_ = ~new_n_n2096_;
  assign new_n_n404_ = ~new_n_n2472_;
  assign new_n_n394_ = ~new_n_n2110_;
  assign new_n_n384_ = ~new_n_n1625_;
  assign new_n_n374_ = ~new_n_n1626_;
  assign new_n_n350_ = ~new_n_n2145_;
  assign new_n_n340_ = ~new_n_n1621_;
  assign new_n_n331_ = ~new_n_n2152_;
  assign new_n_n323_ = ~new_n_n2163_;
  assign new_n_n320_ = ~new_n_n1615_;
  assign new_n_n310_ = ~new_n_n2175_;
  assign new_n_n300_ = ~new_nb10_;
  assign new_n_n290_ = ~new_n_n2194_;
  assign new_n_n275_ = ~new_n_n2209_;
  assign new_n_n262_ = ~new_n_n2224_;
  assign new_n_n252_ = ~new_n_n2229_;
  assign new_n_n242_ = ~new_n_n2242_;
  assign new_n_n231_ = ~new_n_n1608_;
  assign new_n_n218_ = ~new_n_n1607_;
  assign new_n_n208_ = ~new_n_n2272_;
  assign new_n_n197_ = ~new_n_n2282_;
  assign new_n_n182_ = ~new_n_n1605_;
  assign new_n_n172_ = ~new_n_n2306_;
  assign new_n_n169_ = ~new_n_n1604_;
  assign new_n_n159_ = ~new_n_n2318_;
  assign new_n_n149_ = ~new_n_n2330_;
  assign new_n_n139_ = ~new_n_n2338_;
  assign new_n_n116_ = ~new_nina14_;
  assign new_n_n105_ = ~new_nb15_;
  assign new_n_n1_ = ~new_n_n2486_;
  assign new_n_n2478_ = new_n_n1593_ | new_n_n1594_;
  assign new_n_n2472_ = new_n_n1591_ | new_n_n10_;
  assign new_n_n1588_ = new_n_n18_ & new_n_n1714_;
  assign new_n_n2433_ = new_n_n1714_ | new_n_n815_ | new_n_n295_;
  assign new_n_n2426_ = new_n_n1576_ | new_n_n47_;
  assign new_n_n1573_ = new_n_n56_ & new_n_n840_;
  assign new_n_n1571_ = new_n_n61_ & new_n_n840_;
  assign new_n_n2406_ = new_n_n64_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2399_ = new_n_n840_ | new_n_n71_;
  assign new_n_n2390_ = new_n_n1641_ | new_n_n404_ | new_n_n1642_ | new_n_n366_;
  assign new_n_n2383_ = new_n_n351_ & new_n_n853_ & new_n_n86_;
  assign new_n_n1549_ = new_n_n97_ & new_n_n98_;
  assign new_n_n1547_ = new_n_n104_ & new_n_n105_;
  assign new_n_n1544_ = new_n_n116_ & new_n_n1714_;
  assign new_n_n2358_ = new_n_n1715_ | new_n_n820_ | new_n_n357_;
  assign new_n_n2352_ = new_n_n123_ & new_n_n815_;
  assign new_n_n2350_ = new_n_n125_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n1522_ = new_n_n142_ & new_n_n1714_;
  assign new_n_n2334_ = new_n_n815_ | new_n_n1713_ | new_n_n1634_;
  assign new_n_n1510_ = new_n_n157_ & new_n_n1715_;
  assign new_n_n1506_ = new_n_n153_ & new_n_n154_;
  assign new_n_n1505_ = new_n_n79_ & new_n_n158_;
  assign new_n_n1500_ = new_n_n815_ & new_n_n1604_;
  assign new_n_n2307_ = new_n_n169_ & new_n_n815_;
  assign new_n_n1490_ = new_n_n104_ & new_n_n175_;
  assign new_n_n1470_ = new_n_n1714_ & new_n_n191_;
  assign new_n_n1465_ = new_n_n2159_ & new_nb0_;
  assign new_n_n2275_ = new_n_n1712_ & new_n_n801_;
  assign new_n_n2260_ = new_n_n218_ & new_n_n815_;
  assign new_n_n1418_ = new_n_n2159_ & new_nb5_;
  assign new_n_n2227_ = new_n_n1412_ | new_n_n1413_;
  assign new_n_n2021_ = new_n_n500_ | new_n_n501_;
  assign new_n_n2016_ = new_n_n1180_ | new_n_n1181_;
  assign new_n_n1986_ = new_n_n1724_ | new_n_n539_;
  assign new_n_n1975_ = new_n_n1659_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1135_ = new_n_n533_ & new_n_n557_;
  assign new_n_n1964_ = new_n_n1126_ | new_n_n1127_;
  assign new_n_n1121_ = new_n_n568_ & new_n_n571_;
  assign new_n_n1948_ = new_n_n1103_ | new_n_n879_ | new_n_n1104_ | new_n_n1105_;
  assign new_n_n1100_ = new_n_n836_ & new_n_n589_;
  assign new_n_n1094_ = new_n_n596_ & new_n_n351_;
  assign new_n_n1933_ = new_n_n1088_ | new_n_n1089_;
  assign new_n_n1087_ = new_n_n603_ & new_n_n604_;
  assign new_n_n1082_ = new_n_n612_ & new_n_n611_;
  assign new_n_n1075_ = new_n_n621_ & new_n_n1714_;
  assign new_n_n1071_ = new_n_n831_ & new_n_n716_;
  assign new_n_n1906_ = new_n_n675_ | new_n_n1684_;
  assign new_n_n1901_ = new_n_n1056_ | new_n_n1057_;
  assign new_n_n1053_ = new_n_n649_ & new_n_n648_;
  assign new_n_n1893_ = new_n_n1680_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1042_ = new_n_n833_ & new_n_n662_;
  assign new_n_n1039_ = new_n_n833_ & new_n_n664_;
  assign new_n_n1028_ = new_n_n1734_ & new_n_n1684_;
  assign new_n_n1872_ = new_n_n1021_ | new_n_n1022_;
  assign new_n_n1015_ = new_n_n756_ & new_n_n1719_;
  assign new_n_n1010_ = new_n_n833_ & new_n_n691_;
  assign new_n_n1859_ = new_n_n1005_ | new_n_n1006_;
  assign new_n_n1000_ = new_n_n568_ & new_n_n702_;
  assign new_n_n992_ = new_n_n705_ & new_n_n706_;
  assign new_n_n1849_ = new_n_n1694_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1822_ = new_n_n747_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n1818_ = new_n_n958_ | new_n_n753_;
  assign new_n_n1805_ = new_n_n767_ & new_n_n351_;
  assign new_n_n911_ = new_n_n796_ & new_n_n1724_;
  assign new_n_n1773_ = new_n_n907_ | new_n_n908_;
  assign new_n_n816_ = ~new_n_n1714_;
  assign new_n_n807_ = ~new_n_n1771_;
  assign new_n_n797_ = ~new_n_n1779_;
  assign new_n_n789_ = ~new_n_n1786_;
  assign new_n_n755_ = ~new_n_n1817_;
  assign new_n_n730_ = ~new_n_n1802_;
  assign new_n_n724_ = ~new_n_n1838_;
  assign new_n_n713_ = ~new_n_n1850_;
  assign new_n_n705_ = ~new_n_n1853_;
  assign new_n_n682_ = ~new_n_n1878_;
  assign new_n_n1683_ = ~new_n_n1885_;
  assign new_n_n651_ = ~new_n_n1676_;
  assign new_n_n643_ = ~new_n_n1678_;
  assign new_n_n634_ = ~new_n_n2454_;
  assign new_n_n626_ = ~new_n_n1919_;
  assign new_n_n1670_ = ~new_n_n2263_;
  assign new_n_n592_ = ~new_n_n1944_;
  assign new_n_n572_ = ~new_n_n1960_;
  assign new_n_n570_ = ~new_n_n1663_;
  assign new_n_n562_ = ~new_n_n1966_;
  assign new_n_n551_ = ~new_n_n1659_;
  assign new_n_n1658_ = ~new_n_n2179_;
  assign new_n_n516_ = ~new_n_n2006_;
  assign new_n_n507_ = ~new_n_n2011_;
  assign new_n_n496_ = ~new_n_n1995_;
  assign new_n_n1648_ = ~new_nind10_;
  assign new_n_n485_ = ~new_n_n2033_;
  assign new_n_n476_ = ~new_n_n2037_;
  assign new_n_n1646_ = ~new_n_n2057_;
  assign new_n_n457_ = ~new_n_n2056_;
  assign new_n_n1639_ = ~new_n_n2077_;
  assign new_n_n424_ = ~new_n_n2063_;
  assign new_n_n414_ = ~new_n_n2088_;
  assign new_n_n407_ = ~new_n_n2095_;
  assign new_n_n403_ = ~new_n_n2100_;
  assign new_n_n395_ = ~new_n_n2106_;
  assign new_n_n383_ = ~new_n_n2118_;
  assign new_n_n375_ = ~new_n_n1627_;
  assign new_n_n349_ = ~new_n_n2141_;
  assign new_n_n341_ = ~new_n_n1740_;
  assign new_n_n1618_ = ~new_n_n2186_;
  assign new_n_n324_ = ~new_n_n2162_;
  assign new_n_n1615_ = ~new_ninc8_;
  assign new_n_n311_ = ~new_n_n2174_;
  assign new_n_n299_ = ~new_n_n2190_;
  assign new_n_n291_ = ~new_n_n2193_;
  assign new_n_n266_ = ~new_n_n1906_;
  assign new_n_n261_ = ~new_n_n2221_;
  assign new_n_n253_ = ~new_n_n2228_;
  assign new_n_n241_ = ~new_n_n2239_;
  assign new_n_n232_ = ~new_nina6_;
  assign new_n_n228_ = ~new_n_n2252_;
  assign new_n_n207_ = ~new_n_n2271_;
  assign new_n_n198_ = ~new_n_n2281_;
  assign new_n_n1605_ = ~new_ninc1_;
  assign new_n_n173_ = ~new_n_n2305_;
  assign new_n_n1604_ = ~new_ninc2_;
  assign new_n_n160_ = ~new_n_n2317_;
  assign new_n_n148_ = ~new_n_n2329_;
  assign new_n_n140_ = ~new_n_n2341_;
  assign new_n_n115_ = ~new_nb14_;
  assign new_n_n106_ = ~new_n_n2369_;
  assign new_n_n2_ = ~new_n_n2484_;
  assign new_n_n1594_ = new_n_n1731_ & new_n_n6_;
  assign new_n_n2470_ = new_n_n1714_ | new_n_n815_ | new_n_n142_;
  assign new_n_n2465_ = new_n_n1607_ | new_n_n1715_;
  assign new_n_n2432_ = new_n_n1578_ | new_n_n42_;
  assign new_n_n2424_ = new_n_n840_ | new_n_n51_;
  assign new_n_n2419_ = new_n_n54_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2410_ = new_n_n1571_ | new_n_n60_;
  assign new_n_n2405_ = new_n_n840_ | new_n_n66_;
  assign new_n_n2397_ = new_n_n1606_ | new_n_n1715_;
  assign new_n_n1565_ = new_n_n76_ & new_n_n840_;
  assign new_n_n2378_ = new_n_n1715_ | new_n_n820_ | new_n_n90_;
  assign new_n_n1550_ = new_n_n97_ & new_n_n1714_;
  assign new_n_n2369_ = new_n_n107_ | new_n_n108_;
  assign new_nb14_ = new_n_n113_ & new_n_n114_;
  assign new_n_n1538_ = new_n_n116_ & new_n_n1600_;
  assign new_n_n2353_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n122_;
  assign new_nb13_ = new_n_n126_ & new_n_n127_;
  assign new_n_n2344_ = new_n_n1525_ | new_n_n1526_;
  assign new_n_n1515_ = new_n_n1714_ & new_n_n144_;
  assign new_n_n1512_ = new_n_n148_ & new_n_n149_;
  assign new_n_n2322_ = new_n_n1506_ | new_n_n819_;
  assign new_n_n1504_ = new_n_n157_ & new_n_n1714_;
  assign new_n_n2314_ = new_n_n163_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n1495_ = new_n_n166_ & new_n_n167_;
  assign new_n_n1491_ = new_n_n2159_ & new_nb2_;
  assign new_n_n2284_ = new_n_n1606_ | new_n_n1716_;
  assign new_n_n2280_ = new_n_n198_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2276_ = new_n_n1726_ & new_n_n845_;
  assign new_n_n2267_ = new_n_n212_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2237_ = new_n_n1609_ | new_n_n1716_;
  assign new_n_n2009_ = new_n_n508_ | new_n_n515_;
  assign new_n_n1174_ = new_n_n519_ & new_n_n520_;
  assign new_n_n1980_ = new_n_n1147_ | new_n_n1148_;
  assign new_n_n1974_ = new_n_n1138_ | new_n_n554_;
  assign new_n_n1133_ = new_n_n831_ & new_n_n586_;
  assign new_n_n1966_ = new_n_n563_ | new_n_n564_;
  assign new_n_n1122_ = new_n_n567_ & new_n_n434_;
  assign new_n_n1105_ = new_n_n833_ & new_n_n585_;
  assign new_n_n1943_ = new_n_n592_ | new_n_n593_;
  assign new_n_n1940_ = new_n_n1724_ | new_n_n594_;
  assign new_n_n1090_ = new_n_n1690_ & new_n_n605_;
  assign new_n_n1930_ = new_n_n1085_ | new_n_n1086_;
  assign new_n_n1080_ = new_n_n613_ & new_n_n614_;
  assign new_n_n1924_ = new_n_n620_ & new_n_n815_;
  assign new_n_n1918_ = new_n_n1071_ | new_n_n1015_;
  assign new_n_n1912_ = new_n_n633_ | new_n_n634_;
  assign new_n_n1058_ = new_n_n637_ & new_n_n638_;
  assign new_n_n1057_ = new_n_n1677_ & new_n_n1678_;
  assign new_n_n1051_ = new_n_n351_ & new_n_n651_;
  assign new_n_n1048_ = new_n_n79_ & new_n_n658_;
  assign new_n_n1888_ = new_n_n1040_ | new_n_n879_ | new_n_n1041_ | new_n_n1042_;
  assign new_n_n1038_ = new_n_n665_ & new_n_n664_;
  assign new_n_n1032_ = new_n_n671_ & new_n_n1724_;
  assign new_n_n1023_ = new_n_n676_ & new_n_n677_;
  assign new_n_n1016_ = new_n_n83_ & new_n_n687_;
  assign new_n_n1861_ = new_n_n981_ | new_n_n879_ | new_n_n1009_ | new_n_n1010_;
  assign new_n_n1006_ = new_n_n695_ & new_n_n696_;
  assign new_n_n998_ = new_n_n1691_ & new_n_n700_;
  assign new_n_n1853_ = new_n_n704_ & new_n_n351_;
  assign new_n_n987_ = new_n_n710_ & new_n_n711_;
  assign new_n_n1823_ = new_n_n963_ | new_n_n964_;
  assign new_n_n1819_ = new_n_n1701_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n949_ = new_n_n762_ & new_n_n1721_;
  assign new_n_n815_ = ~new_n_n1715_;
  assign new_n_n804_ = ~new_n_n1727_;
  assign new_n_n1710_ = ~new_n_n1784_;
  assign new_n_n790_ = ~new_n_n1757_;
  assign new_n_n746_ = ~new_ne3_;
  assign new_n_n729_ = ~new_n_n1699_;
  assign new_n_n722_ = ~new_n_n1840_;
  assign new_n_n716_ = ~new_n_n1649_;
  assign new_n_n706_ = ~new_n_n1693_;
  assign new_n_n666_ = ~new_n_n1888_;
  assign new_n_n657_ = ~new_ninb5_;
  assign new_n_n650_ = ~new_n_n1901_;
  assign new_n_n1677_ = ~new_n_n2245_;
  assign new_n_n636_ = ~new_n_n1909_;
  assign new_n_n627_ = ~new_n_n1623_;
  assign new_n_n1669_ = ~new_n_n2257_;
  assign new_n_n583_ = ~new_n_n1954_;
  assign new_n_n573_ = ~new_n_n1958_;
  assign new_n_n569_ = ~new_n_n1662_;
  assign new_n_n559_ = ~new_n_n1949_;
  assign new_n_n1659_ = ~new_nind8_;
  assign new_n_n543_ = ~new_n_n1735_;
  assign new_n_n515_ = ~new_n_n2015_;
  assign new_n_n505_ = ~new_n_n1651_;
  assign new_n_n499_ = ~new_n_n2021_;
  assign new_n_n490_ = ~new_n_n2030_;
  assign new_n_n484_ = ~new_n_n2034_;
  assign new_n_n473_ = ~new_n_n2038_;
  assign new_n_n467_ = ~new_n_n1619_;
  assign new_n_n458_ = ~new_n_n2053_;
  assign new_n_n443_ = ~new_n_n2070_;
  assign new_n_n1638_ = ~new_n_n2331_;
  assign new_n_n422_ = ~new_n_n424_;
  assign new_n_n417_ = ~new_n_n1634_;
  assign new_n_n408_ = ~new_n_n1631_;
  assign new_n_n402_ = ~new_n_n2099_;
  assign new_n_n1629_ = ~new_nind13_;
  assign new_n_n386_ = ~new_ne14_;
  assign new_n_n376_ = ~new_n_n2121_;
  assign new_n_n364_ = ~new_n_n2129_;
  assign new_n_n355_ = ~new_n_n2382_;
  assign new_n_n348_ = ~new_n_n2368_;
  assign new_n_n338_ = ~new_n_n2148_;
  assign new_n_n333_ = ~new_n_n2151_;
  assign new_n_n325_ = ~new_n_n2165_;
  assign new_n_n319_ = ~new_n_n2166_;
  assign new_n_n308_ = ~new_nina9_;
  assign new_n_n302_ = ~new_n_n2182_;
  assign new_n_n292_ = ~new_n_n2196_;
  assign new_n_n277_ = ~new_n_n2206_;
  assign new_n_n267_ = ~new_n_n2216_;
  assign new_n_n260_ = ~new_n_n2222_;
  assign new_n_n250_ = ~new_nb5_;
  assign new_n_n1609_ = ~new_ninc5_;
  assign new_n_n233_ = ~new_n_n2248_;
  assign new_n_n227_ = ~new_n_n2253_;
  assign new_n_n217_ = ~new_n_n2262_;
  assign new_n_n199_ = ~new_n_n2280_;
  assign new_n_n184_ = ~new_n_n2294_;
  assign new_n_n174_ = ~new_n_n2308_;
  assign new_n_n168_ = ~new_n_n2309_;
  assign new_n_n157_ = ~new_nina3_;
  assign new_n_n151_ = ~new_n_n2325_;
  assign new_n_n141_ = ~new_nb12_;
  assign new_n_n134_ = ~new_n_n2347_;
  assign new_n_n124_ = ~new_n_n2352_;
  assign new_n_n3_ = ~new_n_n2481_;
  assign new_n_n1596_ = new_n_n1_ & new_n_n1714_;
  assign new_n_n1593_ = new_n_n1597_ & new_n_n840_;
  assign new_n_n2471_ = new_n_n1602_ | new_n_n1715_;
  assign new_n_n2464_ = new_n_n1714_ | new_n_n815_ | new_n_n219_;
  assign new_n_n1578_ = new_n_n43_ & new_n_n1714_;
  assign new_n_n2425_ = new_n_n49_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2418_ = new_n_n840_ | new_n_n56_;
  assign new_n_n2411_ = new_n_n840_ | new_n_n61_;
  assign new_n_n2404_ = new_n_n1569_ | new_n_n65_;
  assign new_n_n1567_ = new_n_n71_ & new_n_n840_;
  assign new_n_n2391_ = new_n_n1722_ | new_n_n765_ | new_n_n795_ | new_n_n723_;
  assign new_n_n1559_ = new_n_n87_ & new_n_n351_;
  assign new_n_n2377_ = new_n_n1553_ | new_n_n1554_;
  assign new_n_n1551_ = new_n_n79_ & new_n_n98_;
  assign new_n_n2368_ = new_n_n1546_ | new_n_n106_;
  assign new_n_n2363_ = new_n_n112_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2360_ = new_n_n117_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2354_ = new_n_n1601_ | new_n_n1716_;
  assign new_n_n2349_ = new_n_n1530_ | new_n_n1531_;
  assign new_n_n2345_ = new_n_n1715_ | new_n_n820_ | new_n_n391_;
  assign new_n_n2339_ = new_n_n1521_ | new_n_n1523_ | new_n_n1522_ | new_n_n893_;
  assign new_n_n2332_ = new_n_n1514_ | new_n_n1515_;
  assign new_n_n2327_ = new_n_n1509_ | new_n_n1511_ | new_n_n1510_ | new_n_n1358_;
  assign new_n_n1507_ = new_n_n1714_ & new_n_n152_;
  assign new_n_n1503_ = new_n_n157_ & new_n_n158_;
  assign new_n_n1498_ = new_n_n170_ & new_n_n1604_;
  assign new_n_n2309_ = new_n_n1604_ | new_n_n1716_;
  assign new_n_n2304_ = new_n_n1490_ | new_n_n1491_;
  assign new_n_n1469_ = new_n_n192_ & new_n_n193_;
  assign new_nb0_ = new_n_n199_ & new_n_n200_;
  assign new_n_n2277_ = new_n_n203_ | new_n_n202_;
  assign new_n_n2272_ = new_n_n1706_ & new_n_n770_;
  assign new_n_n1422_ = new_n_n241_ & new_n_n242_;
  assign new_n_n2008_ = new_n_n510_ | new_n_n511_;
  assign new_n_n1175_ = new_n_n519_ & new_n_n518_;
  assign new_no9_ = new_n_n1142_ | new_n_n549_;
  assign new_n_n1138_ = new_n_n83_ & new_n_n555_;
  assign new_n_n1969_ = new_n_n1133_ | new_n_n1107_;
  assign new_n_n1965_ = new_n_n1128_ | new_n_n562_;
  assign new_n_n1123_ = new_n_n567_ & new_n_n571_;
  assign new_n_n1104_ = new_n_n559_ & new_n_n585_;
  assign new_n_n1944_ = new_n_n1691_ | new_n_n670_ | new_n_n1692_ | new_n_n634_;
  assign new_n_n1939_ = new_n_n595_ & new_n_n351_;
  assign new_n_n1934_ = new_n_n1090_ | new_n_n644_;
  assign new_n_n1086_ = new_n_n605_ & new_n_n1690_;
  assign new_n_n1081_ = new_n_n613_ & new_n_n612_;
  assign new_n_n1923_ = new_n_n1074_ | new_n_n1076_ | new_n_n1075_ | new_n_n893_;
  assign new_n_n1072_ = new_n_n788_ & new_n_n1719_;
  assign new_n_n1911_ = new_n_n1063_ | new_n_n632_;
  assign new_n_n1059_ = new_n_n637_ & new_n_n351_;
  assign new_n_n1056_ = new_n_n642_ & new_n_n643_;
  assign new_n_n1897_ = new_n_n1050_ | new_n_n1051_;
  assign new_n_n1047_ = new_n_n657_ & new_n_n1714_;
  assign new_n_n1043_ = new_n_n831_ & new_n_n758_;
  assign new_n_n1885_ = new_n_n1036_ | new_n_n1037_;
  assign new_n_n1033_ = new_n_n671_ & new_n_n1683_;
  assign new_n_n1029_ = new_n_n1690_ & new_n_n639_;
  assign new_n_n1866_ = new_n_n1719_ | new_n_n1686_;
  assign new_n_n1862_ = new_n_n1106_ | new_n_n985_;
  assign new_n_n1005_ = new_n_n1687_ & new_n_n1688_;
  assign new_n_n1856_ = new_n_n997_ | new_n_n998_;
  assign new_n_n1852_ = new_n_n992_ | new_n_n993_;
  assign new_n_n988_ = new_n_n710_ & new_n_n1714_;
  assign new_n_n964_ = new_n_n351_ & new_n_n745_;
  assign new_n_n959_ = new_n_n751_ & new_n_n752_;
  assign new_n_n1814_ = new_n_n953_ | new_n_n879_ | new_n_n954_ | new_n_n955_;
  assign new_n_n814_ = ~new_n_n1717_;
  assign new_n_n805_ = ~new_n_n1772_;
  assign new_n_n799_ = ~new_n_n1709_;
  assign new_n_n791_ = ~new_n_n1787_;
  assign new_n_n1700_ = ~new_n_n1803_;
  assign new_n_n728_ = ~new_n_n1698_;
  assign new_n_n723_ = ~new_n_n2410_;
  assign new_n_n715_ = ~new_n_n1846_;
  assign new_n_n707_ = ~new_n_n1857_;
  assign new_n_n665_ = ~new_n_n1864_;
  assign new_n_n658_ = ~new_n_n1895_;
  assign new_n_n649_ = ~new_n_n1898_;
  assign new_n_n1678_ = ~new_n_n2251_;
  assign new_n_n635_ = ~new_n_n1911_;
  assign new_n_n1674_ = ~new_n_n1921_;
  assign new_n_n590_ = ~new_n_n1946_;
  assign new_n_n582_ = ~new_n_n1953_;
  assign new_n_n574_ = ~new_n_n1957_;
  assign new_n_n568_ = ~new_n_n1963_;
  assign new_n_n560_ = ~new_n_n1970_;
  assign new_n_n553_ = ~new_n_n1977_;
  assign new_n_n544_ = ~new_n_n1980_;
  assign new_n_n514_ = ~new_n_n1981_;
  assign new_n_n1652_ = ~new_n_n2023_;
  assign new_n_n498_ = ~new_n_n2024_;
  assign new_n_n491_ = ~new_n_n2031_;
  assign new_n_n483_ = ~new_ne11_;
  assign new_n_n474_ = ~new_n_n1736_;
  assign new_n_n466_ = ~new_n_n1620_;
  assign new_n_n459_ = ~new_n_n2054_;
  assign new_n_n435_ = ~new_n_n1642_;
  assign new_n_n1637_ = ~new_n_n2337_;
  assign new_n_n1636_ = ~new_n_n2083_;
  assign new_n_n416_ = ~new_n_n2094_;
  assign new_n_n1632_ = ~new_n_n2101_;
  assign new_n_n401_ = ~new_n_n2112_;
  assign new_n_n393_ = ~new_n_n2109_;
  assign new_n_n385_ = ~new_n_n1770_;
  assign new_n_n1628_ = ~new_n_n2093_;
  assign new_n_n363_ = ~new_n_n2133_;
  assign new_n_n356_ = ~new_n_n1622_;
  assign new_n_n347_ = ~new_n_n2142_;
  assign new_n_n339_ = ~new_n_n2147_;
  assign new_n_n332_ = ~new_n_n2153_;
  assign new_n_n326_ = ~new_n_n1730_;
  assign new_n_n318_ = ~new_n_n2171_;
  assign new_n_n309_ = ~new_n_n2176_;
  assign new_n_n301_ = ~new_n_n2184_;
  assign new_n_n293_ = ~new_n_n2191_;
  assign new_n_n276_ = ~new_n_n2207_;
  assign new_n_n268_ = ~new_n_n2217_;
  assign new_n_n259_ = ~new_n_n2223_;
  assign new_n_n251_ = ~new_n_n2231_;
  assign new_n_n243_ = ~new_n_n2237_;
  assign new_n_n234_ = ~new_n_n2247_;
  assign new_n_n226_ = ~new_n_n2254_;
  assign new_n_n1607_ = ~new_ninc7_;
  assign new_n_n209_ = ~new_n_n2273_;
  assign new_n_n183_ = ~new_nina1_;
  assign new_n_n175_ = ~new_nb2_;
  assign new_n_n167_ = ~new_n_n2314_;
  assign new_n_n158_ = ~new_n_n2319_;
  assign new_n_n150_ = ~new_n_n2327_;
  assign new_n_n142_ = ~new_nina12_;
  assign new_n_n133_ = ~new_n_n2344_;
  assign new_n_n125_ = ~new_n_n2351_;
  assign new_n_n4_ = ~new_n_n2482_;
  assign new_n_n2482_ = new_n_n1599_ | new_n_n1715_;
  assign new_n_n1592_ = new_n_n8_ & new_n_n1714_;
  assign new_n_n2466_ = new_n_n1589_ | new_n_n15_;
  assign new_n_n2393_ = new_n_n840_ | new_n_n76_;
  assign new_n_n1372_ = new_n_n1647_ & new_n_n466_;
  assign new_n_n1366_ = new_n_n1714_ & new_n_n302_;
  assign new_n_n2174_ = new_n_n310_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n1323_ = new_n_n349_ & new_n_n348_;
  assign new_n_n1317_ = new_n_n357_ & new_n_n1714_;
  assign new_n_n2132_ = new_n_n363_ | new_n_n1635_;
  assign new_n_n2126_ = new_n_n1724_ | new_n_n367_;
  assign new_n_n1303_ = new_n_n1626_ & new_n_n1627_;
  assign new_n_n1297_ = new_n_n351_ & new_n_n384_;
  assign new_n_n2093_ = new_n_n2331_ | new_n_n1637_;
  assign new_n_n1271_ = new_n_n410_ & new_n_n372_;
  assign new_n_n1265_ = new_n_n418_ & new_n_n1714_;
  assign new_n_n1258_ = new_n_n690_ & new_n_n1720_;
  assign new_n_n2077_ = new_n_n1249_ | new_n_n1250_;
  assign new_n_n1243_ = new_n_n1641_ & new_n_n435_;
  assign new_no12_ = new_n_n1235_ | new_n_n1236_;
  assign new_n_n2065_ = new_n_n627_ & new_n_n1719_;
  assign new_n_n1226_ = new_n_n423_ & new_n_n690_;
  assign new_n_n1211_ = new_n_n469_ & new_n_n274_;
  assign new_n_n2037_ = new_n_n1205_ | new_n_n472_;
  assign new_n_n1199_ = new_n_n385_ & new_n_n483_;
  assign new_n_n1194_ = new_n_n83_ & new_n_n491_;
  assign new_n_n1188_ = new_n_n496_ & new_n_n495_;
  assign new_n_n1182_ = new_n_n502_ & new_n_n1724_;
  assign new_n_n1179_ = new_n_n1616_ & new_n_n506_;
  assign new_ne10_ = new_n_n1174_ | new_n_n1175_;
  assign new_n_n1148_ = new_n_n545_ & new_n_n513_;
  assign new_n_n1977_ = new_n_n551_ & new_n_n815_;
  assign new_n_n1137_ = new_n_n831_ & new_n_n663_;
  assign new_n_n1130_ = new_n_n836_ & new_n_n560_;
  assign new_n_n1962_ = new_n_n999_ | new_n_n1122_ | new_n_n1121_ | new_n_n1123_;
  assign new_no7_ = new_n_n1077_ | new_n_n618_;
  assign new_n_n1919_ = new_n_n1072_ | new_n_n625_;
  assign new_n_n92_ = ~new_n_n2378_;
  assign new_n_n82_ = ~new_n_n2387_;
  assign new_n_n71_ = ~new_n_n2400_;
  assign new_n_n60_ = ~new_n_n2411_;
  assign new_n_n49_ = ~new_n_n2426_;
  assign new_n_n2481_ = new_n_n1714_ | new_n_n815_ | new_n_n97_;
  assign new_n_n2475_ = new_n_n1592_ | new_n_n7_;
  assign new_n_n1589_ = new_n_n16_ & new_n_n840_;
  assign new_n_n2392_ = new_n_n1565_ | new_n_n75_;
  assign new_n_n1371_ = new_n_n510_ & new_n_n1619_;
  assign new_n_n2180_ = new_n_n1365_ | new_n_n1366_;
  assign new_n_n2171_ = new_n_n314_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n1322_ = new_n_n349_ & new_n_n350_;
  assign new_n_n1318_ = new_n_n79_ & new_n_n358_;
  assign new_n_n2131_ = new_n_n1310_ | new_n_n362_;
  assign new_n_n1306_ = new_n_n367_ & new_n_n1724_;
  assign new_n_n1302_ = new_n_n374_ & new_n_n375_;
  assign new_n_n2114_ = new_n_n1296_ | new_n_n1297_;
  assign new_n_n2092_ = new_n_n1276_ | new_n_n376_;
  assign new_ne13_ = new_n_n1270_ | new_n_n1271_;
  assign new_n_n1264_ = new_n_n418_ & new_n_n419_;
  assign new_n_n2081_ = new_n_n1257_ | new_n_n1258_;
  assign new_n_n1250_ = new_n_n429_ & new_n_n430_;
  assign new_n_n2074_ = new_n_n1242_ | new_n_n1243_;
  assign new_n_n1236_ = new_n_n576_ & new_n_n442_;
  assign new_n_n1231_ = new_n_n83_ & new_n_n448_;
  assign new_n_n2055_ = new_n_n457_ | new_n_n840_;
  assign new_n_n2042_ = new_n_n1209_ | new_n_n1210_;
  assign new_n_n1206_ = new_n_n506_ & new_n_n512_;
  assign new_n_n2033_ = new_n_n484_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n2029_ = new_n_n1194_ | new_n_n490_;
  assign new_n_n2023_ = new_n_n1186_ | new_n_n1187_;
  assign new_n_n1183_ = new_n_n502_ & new_n_n1652_;
  assign new_n_n2010_ = new_n_n507_ | new_n_n472_;
  assign new_n_n1176_ = new_n_n520_ & new_n_n517_;
  assign new_n_n1985_ = new_n_n540_ & new_n_n351_;
  assign new_n_n1976_ = new_n_n1139_ | new_n_n1141_ | new_n_n1140_ | new_n_n893_;
  assign new_n_n1971_ = new_n_n1137_ | new_n_n1072_;
  assign new_n_n1129_ = new_n_n561_ & new_n_n1721_;
  assign new_n_n1124_ = new_n_n849_ & new_n_n1729_;
  assign new_n_n1077_ = new_n_n619_ & new_n_n1730_;
  assign new_n_n1920_ = new_n_n1719_ | new_n_n1674_;
  assign new_n_n93_ = ~new_n_n2377_;
  assign new_n_n81_ = ~new_n_n1762_;
  assign new_n_n72_ = ~new_n_n2396_;
  assign new_n_n59_ = ~new_n_n2413_;
  assign new_n_n50_ = ~new_n_n2424_;
  assign new_n_n2480_ = new_n_n1595_ | new_n_n3_;
  assign new_n_n2473_ = new_n_n840_ | new_n_n11_;
  assign new_n_n2468_ = new_n_n14_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2408_ = new_n_n1714_ | new_n_n815_ | new_n_n170_;
  assign new_n_n2400_ = new_n_n69_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2185_ = new_n_n1370_ | new_n_n1372_ | new_n_n1371_ | new_n_n1373_;
  assign new_n_n2181_ = new_n_n1715_ | new_n_n820_ | new_n_n527_;
  assign new_n_n2164_ = new_n_n320_ & new_n_n815_;
  assign new_n_n1324_ = new_n_n348_ & new_n_n347_;
  assign new_n_n2137_ = new_n_n1316_ | new_n_n1318_ | new_n_n1317_ | new_n_n893_;
  assign new_n_n1310_ = new_n_n363_ & new_n_n627_;
  assign new_n_n2124_ = new_n_n1304_ | new_n_n1305_;
  assign new_n_n2119_ = new_n_n373_ | new_n_n378_;
  assign new_n_n1298_ = new_n_n382_ & new_n_n383_;
  assign new_n_n1272_ = new_n_n411_ & new_n_n377_;
  assign new_n_n2084_ = new_n_n1634_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n2080_ = new_n_n1255_ | new_n_n1256_;
  assign new_n_n1252_ = new_n_n831_ & new_n_n427_;
  assign new_n_n1244_ = new_n_n568_ & new_n_n437_;
  assign new_n_n1235_ = new_n_n443_ & new_n_n1730_;
  assign new_n_n1227_ = new_n_n450_ & new_n_n1649_;
  assign new_n_n2056_ = new_n_n856_ & new_n_n456_;
  assign new_n_n1210_ = new_n_n474_ & new_n_n472_;
  assign new_n_n2036_ = new_n_n476_ | new_n_n475_;
  assign new_n_n2034_ = new_n_n1199_ | new_n_n1200_;
  assign new_n_n2030_ = new_n_n1648_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n1187_ = new_n_n836_ & new_n_n497_;
  assign new_n_n2017_ = new_n_n503_ & new_n_n351_;
  assign new_n_n2012_ = new_n_n563_ | new_n_n1657_;
  assign new_n_n1177_ = new_n_n520_ & new_n_n472_;
  assign new_n_n1157_ = new_n_n535_ & new_n_n1721_;
  assign new_n_n1141_ = new_n_n79_ & new_n_n553_;
  assign new_n_n1136_ = new_n_n833_ & new_n_n557_;
  assign new_n_n1131_ = new_n_n559_ & new_n_n558_;
  assign new_n_n1125_ = new_n_n848_ & new_n_n1728_;
  assign new_n_n1088_ = new_n_n608_ & new_n_n602_;
  assign new_n_n1083_ = new_n_n612_ & new_n_n1672_;
  assign new_n_n94_ = ~new_n_n2380_;
  assign new_n_n80_ = ~new_n_n2389_;
  assign new_n_n69_ = ~new_n_n2401_;
  assign new_n_n62_ = ~new_n_n2408_;
  assign new_n_n51_ = ~new_n_n2425_;
  assign new_n_n1595_ = new_n_n4_ & new_n_n1714_;
  assign new_n_n2474_ = new_n_n9_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n2467_ = new_n_n840_ | new_n_n16_;
  assign new_n_n2407_ = new_n_n1570_ | new_n_n62_;
  assign new_n_n1568_ = new_n_n68_ & new_n_n1714_;
  assign new_n_n1373_ = new_n_n1647_ & new_n_n1619_;
  assign new_n_n2182_ = new_n_n815_ | new_n_n1713_ | new_n_n1653_;
  assign new_n_n2160_ = new_n_n853_ & new_n_n326_;
  assign new_ne15_ = new_n_n1322_ | new_n_n1323_;
  assign new_n_n2138_ = new_n_n356_ & new_n_n815_;
  assign new_n_n2130_ = new_n_n1641_ | new_n_n404_ | new_n_n1642_;
  assign new_n_n2125_ = new_n_n368_ & new_n_n351_;
  assign new_n_n2118_ = new_n_n1302_ | new_n_n1303_;
  assign new_n_n1299_ = new_n_n382_ & new_n_n381_;
  assign new_n_n1277_ = new_n_n407_ & new_n_n408_;
  assign new_n_n2083_ = new_n_n1263_ | new_n_n420_;
  assign new_n_n1257_ = new_n_n833_ & new_n_n627_;
  assign new_n_n1251_ = new_n_n428_ & new_n_n1719_;
  assign new_n_n1245_ = new_n_n433_ & new_n_n434_;
  assign new_n_n2064_ = new_n_n1229_ | new_n_n1230_;
  assign new_n_n2059_ = new_n_n1225_ | new_n_n1226_;
  assign new_n_n1220_ = new_n_n424_ & new_n_n455_;
  assign new_n_n1209_ = new_n_n474_ & new_n_n507_;
  assign new_n_n1205_ = new_n_n473_ & new_n_n474_;
  assign new_n_n1200_ = new_n_n351_ & new_n_n482_;
  assign new_n_n1195_ = new_n_n488_ & new_n_n489_;
  assign new_n_n1186_ = new_n_n498_ & new_n_n1721_;
  assign new_n_n2018_ = new_n_n1724_ | new_n_n502_;
  assign new_n_n2011_ = new_n_n1179_ | new_n_n512_;
  assign new_n_n2004_ = new_n_n1176_ | new_n_n1177_;
  assign new_n_n1164_ = new_n_n833_ & new_n_n532_;
  assign new_n_n1140_ = new_n_n552_ & new_n_n1714_;
  assign new_n_n1970_ = new_n_n1134_ | new_n_n879_ | new_n_n1135_ | new_n_n1136_;
  assign new_n_n1967_ = new_n_n1129_ | new_n_n1130_;
  assign new_n_n1963_ = new_n_n1124_ | new_n_n1125_;
  assign new_n_n1932_ = new_n_n642_ | new_n_n1678_;
  assign new_n_n1927_ = new_n_n1082_ | new_n_n1083_;
  assign new_n_n95_ = ~new_n_n2375_;
  assign new_n_n79_ = ~new_n_n1765_;
  assign new_n_n70_ = ~new_n_n2399_;
  assign new_n_n61_ = ~new_n_n2412_;
  assign new_n_n52_ = ~new_n_n2421_;
  assign new_n_n0_ = ~new_n_n2485_;
  assign new_n_n2423_ = new_n_n1575_ | new_n_n50_;
  assign new_n_n2415_ = new_n_n1603_ | new_n_n1715_;
  assign new_n_n1419_ = new_n_n245_ & new_n_n246_;
  assign new_n_n2229_ = new_n_n815_ | new_n_n1713_ | new_n_n1685_;
  assign new_n_n1410_ = new_n_n79_ & new_n_n259_;
  assign new_n_n1375_ = new_n_n2159_ & new_nb10_;
  assign new_n_n2183_ = new_n_n301_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2156_ = new_n_n1616_ | new_n_n328_ | new_n_n329_;
  assign new_n_n2141_ = new_n_n1324_ | new_n_n1325_;
  assign new_n_n1319_ = new_n_n355_ & new_n_n1730_;
  assign new_n_n2110_ = new_n_n1292_ | new_n_n1294_ | new_n_n1293_ | new_n_n893_;
  assign new_n_n2104_ = new_n_n1288_ | new_n_n1289_;
  assign new_n_n2100_ = new_n_n1641_ | new_n_n1642_;
  assign new_n_n1278_ = new_n_n407_ & new_n_n351_;
  assign new_n_n1263_ = new_n_n83_ & new_n_n421_;
  assign new_n_n1255_ = new_n_n424_ & new_n_n586_;
  assign new_n_n1248_ = new_n_n1639_ & new_n_n431_;
  assign new_n_n2071_ = new_n_n439_ & new_n_n351_;
  assign new_n_n1232_ = new_n_n445_ & new_n_n446_;
  assign new_n_n2060_ = new_n_n1227_ | new_n_n1228_;
  assign new_n_n2057_ = new_n_n1220_ | new_n_n454_;
  assign new_n_n2041_ = new_n_n2186_ | new_n_n1647_;
  assign new_n_n1204_ = new_n_n479_ & new_n_n477_;
  assign new_n_n2032_ = new_n_n487_ & new_n_n815_;
  assign new_n_n2026_ = new_n_n1190_ | new_n_n879_ | new_n_n1191_ | new_n_n1192_;
  assign new_n_n1190_ = new_n_n494_ & new_n_n1720_;
  assign new_n_n1185_ = new_n_n500_ & new_n_n501_;
  assign new_n_n2014_ = new_n_n2179_ | new_n_n1735_;
  assign new_n_n2005_ = new_n_n516_ | new_n_n515_;
  assign new_n_n1163_ = new_n_n496_ & new_n_n532_;
  assign new_n_n1989_ = new_n_n537_ | new_n_n538_;
  assign new_n_n1151_ = new_n_n541_ & new_n_n542_;
  assign new_n_n1145_ = new_n_n544_ & new_n_n545_;
  assign new_n_n1126_ = new_n_n1616_ & new_n_n566_;
  assign new_n_n1942_ = new_n_n1098_ | new_n_n591_;
  assign new_n_n1937_ = new_n_n1091_ | new_n_n1092_;
  assign new_n_n1775_ = new_n_n772_ | new_n_n1727_;
  assign new_n_n903_ = new_n_n807_ & new_n_n808_;
  assign new_n_n803_ = ~new_n_n1776_;
  assign new_n_n1709_ = ~new_n_n1780_;
  assign new_n_n1694_ = ~new_nind3_;
  assign new_n_n1599_ = ~new_ninc15_;
  assign new_n_n42_ = ~new_n_n2433_;
  assign new_n_n31_ = ~new_n_n2450_;
  assign new_n_n20_ = ~new_n_n2461_;
  assign new_n_n9_ = ~new_n_n2475_;
  assign new_n_n1590_ = new_n_n13_ & new_n_n1714_;
  assign new_n_n1575_ = new_n_n51_ & new_n_n840_;
  assign new_n_n2416_ = new_n_n1663_ | new_n_n501_ | new_n_n538_ | new_n_n460_;
  assign new_n_n1467_ = new_n_n196_ & new_n_n1714_;
  assign new_n_n1420_ = new_n_n245_ & new_n_n1714_;
  assign new_n_n2228_ = new_n_n1715_ | new_n_n820_ | new_n_n684_;
  assign new_n_n2222_ = new_n_n1408_ | new_n_n1410_ | new_n_n1409_ | new_n_n893_;
  assign new_n_n1374_ = new_n_n104_ & new_n_n300_;
  assign new_n_n1367_ = new_n_n308_ & new_n_n1614_;
  assign new_n_n2150_ = new_n_n1212_ | new_n_n333_;
  assign new_n_n1325_ = new_n_n348_ & new_n_n1621_;
  assign new_no15_ = new_n_n1319_ | new_n_n354_;
  assign new_n_n1294_ = new_n_n79_ & new_n_n392_;
  assign new_n_n1290_ = new_n_n831_ & new_n_n1720_;
  assign new_n_n2099_ = new_n_n403_ | new_n_n404_;
  assign new_n_n2094_ = new_n_n1277_ | new_n_n1278_;
  assign new_n_n2082_ = new_n_n1259_ | new_n_n1261_ | new_n_n1260_ | new_n_n1262_;
  assign new_n_n1256_ = new_n_n423_ & new_n_n663_;
  assign new_n_n1241_ = new_n_n853_ & new_n_n437_;
  assign new_n_n2070_ = new_n_n1237_ | new_n_n1238_;
  assign new_n_n1233_ = new_n_n445_ & new_n_n1714_;
  assign new_n_n1228_ = new_n_n450_ & new_n_n833_;
  assign new_n_n1221_ = new_n_n452_ & new_n_n453_;
  assign new_n_n2040_ = new_n_n1208_ | new_n_n475_;
  assign new_n_n2035_ = new_n_n1203_ | new_n_n1204_;
  assign new_n_n2031_ = new_n_n1195_ | new_n_n1197_ | new_n_n1196_ | new_n_n893_;
  assign new_n_n1193_ = new_n_n663_ & new_n_n1719_;
  assign new_n_n2025_ = new_n_n1133_ | new_n_n1166_;
  assign new_n_n2020_ = new_n_n1185_ | new_n_n499_;
  assign new_n_n2013_ = new_n_n1657_ & new_n_n563_;
  assign new_n_n2006_ = new_n_n514_ | new_n_n513_;
  assign new_n_n1162_ = new_n_n496_ & new_n_n1720_;
  assign new_n_n1990_ = new_n_n569_ | new_n_n1663_;
  assign new_n_n1983_ = new_n_n1149_ | new_n_n1150_;
  assign new_n_n1146_ = new_n_n544_ & new_n_n507_;
  assign new_n_n1132_ = new_n_n833_ & new_n_n558_;
  assign new_n_n1098_ = new_n_n592_ & new_n_n593_;
  assign new_n_n1093_ = new_n_n596_ & new_n_n597_;
  assign new_n_n1774_ = new_n_n800_ | new_n_n803_;
  assign new_n_n904_ = new_n_n807_ & new_n_n806_;
  assign new_n_n802_ = ~new_n_n1712_;
  assign new_n_n796_ = ~new_n_n1781_;
  assign new_n_n720_ = ~new_n_n1842_;
  assign new_n_n96_ = ~new_n_n1599_;
  assign new_n_n41_ = ~new_n_n2437_;
  assign new_n_n32_ = ~new_n_n2446_;
  assign new_n_n19_ = ~new_n_n2463_;
  assign new_n_n10_ = ~new_n_n2473_;
  assign new_n_n2476_ = new_n_n1714_ | new_n_n815_ | new_n_n129_;
  assign new_n_n2438_ = new_n_n1580_ | new_n_n37_;
  assign new_n_n2430_ = new_n_n840_ | new_n_n46_;
  assign new_n_n1461_ = new_n_n845_ & new_n_n1712_;
  assign new_nb5_ = new_n_n248_ & new_n_n249_;
  assign new_n_n1414_ = new_n_n258_ & new_n_n1610_;
  assign new_n_n2223_ = new_n_n257_ & new_n_n815_;
  assign new_nb10_ = new_n_n298_ & new_n_n299_;
  assign new_n_n1368_ = new_n_n308_ & new_n_n1715_;
  assign new_n_n1331_ = new_n_n344_ & new_n_n342_;
  assign new_n_n1293_ = new_n_n391_ & new_n_n1714_;
  assign new_n_n1288_ = new_n_n836_ & new_n_n627_;
  assign new_n_n2101_ = new_n_n1283_ | new_n_n399_;
  assign new_n_n2095_ = new_n_n406_ & new_n_n351_;
  assign new_n_n1262_ = new_n_n1635_ & new_n_n1636_;
  assign new_n_n1249_ = new_n_n1637_ & new_n_n1638_;
  assign new_n_n2073_ = new_n_n1239_ | new_n_n913_ | new_n_n1240_ | new_n_n1241_;
  assign new_n_n1238_ = new_n_n440_ & new_n_n351_;
  assign new_n_n2066_ = new_n_n1231_ | new_n_n447_;
  assign new_n_n2062_ = new_n_n1721_ | new_n_n833_;
  assign new_n_n1222_ = new_n_n452_ & new_n_n424_;
  assign new_n_n1208_ = new_n_n470_ & new_n_n471_;
  assign new_ne11_ = new_n_n1201_ | new_n_n1202_;
  assign new_no11_ = new_n_n1198_ | new_n_n485_;
  assign new_n_n2027_ = new_n_n1193_ | new_n_n492_;
  assign new_n_n2024_ = new_n_n1162_ | new_n_n879_ | new_n_n1188_ | new_n_n1189_;
  assign new_n_n1184_ = new_n_n853_ & new_n_n1652_;
  assign new_n_n1180_ = new_n_n504_ & new_n_n505_;
  assign new_n_n1178_ = new_n_n510_ & new_n_n511_;
  assign new_n_n1993_ = new_n_n1133_ | new_n_n1161_;
  assign new_n_n1156_ = new_n_n537_ & new_n_n538_;
  assign new_n_n1984_ = new_n_n1151_ | new_n_n1152_;
  assign new_ne9_ = new_n_n1145_ | new_n_n1146_;
  assign new_n_n1972_ = new_n_n1161_ | new_n_n556_;
  assign new_n_n1952_ = new_n_n1108_ | new_n_n582_;
  assign new_n_n1947_ = new_n_n1133_ | new_n_n1072_;
  assign new_n_n961_ = new_n_n79_ & new_n_n752_;
  assign new_n_n909_ = new_n_n798_ & new_n_n799_;
  assign new_ne1_ = new_n_n903_ | new_n_n904_;
  assign new_n_n820_ = ~new_n_n1713_;
  assign new_n_n812_ = ~new_n_n1768_;
  assign new_n_n1698_ = ~new_n_n2316_;
  assign new_n_n40_ = ~new_n_n2436_;
  assign new_n_n29_ = ~new_n_n2451_;
  assign new_n_n22_ = ~new_n_n2458_;
  assign new_n_n11_ = ~new_n_n2474_;
  assign new_n_n2483_ = new_n_n2_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n1580_ = new_n_n38_ & new_n_n1714_;
  assign new_n_n2431_ = new_n_n44_ | new_n_n820_ | new_n_n1716_;
  assign new_n_n1456_ = new_n_n206_ & new_n_n770_;
  assign new_n_n2233_ = new_n_n247_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2230_ = new_n_n251_ & new_n_n1713_ & new_n_n816_;
  assign new_n_n2224_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n256_;
  assign new_n_n2186_ = new_n_n1374_ | new_n_n1375_;
  assign new_n_n1369_ = new_n_n815_ & new_n_n1614_;
  assign new_n_n2142_ = new_n_n346_ | new_n_n345_;
  assign new_n_n1292_ = new_n_n391_ & new_n_n392_;
  assign new_n_n1289_ = new_n_n663_ & new_n_n1721_;
  assign new_n_n1283_ = new_n_n400_ & new_n_n401_;
  assign new_n_n2096_ = new_n_n1724_ | new_n_n405_;
  assign new_n_n2079_ = new_n_n1253_ | new_n_n1254_;
  assign new_n_n2076_ = new_n_n1247_ | new_n_n1248_;
  assign new_n_n1242_ = new_n_n436_ & new_n_n1642_;
  assign new_n_n1237_ = new_n_n440_ & new_n_n441_;
  assign new_n_n2067_ = new_n_n1644_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n2061_ = new_n_n833_ & new_n_n663_;
  assign new_n_n1223_ = new_n_n831_ & new_n_n453_;
  assign new_n_n2039_ = new_n_n2192_ | new_n_n1618_;
  assign new_n_n1203_ = new_n_n479_ & new_n_n478_;
  assign new_n_n1198_ = new_n_n486_ & new_n_n1730_;
  assign new_n_n2028_ = new_n_n1719_ | new_n_n1650_;
  assign new_n_n1189_ = new_n_n833_ & new_n_n495_;
  assign new_n_n2019_ = new_n_n1182_ | new_n_n913_ | new_n_n1183_ | new_n_n1184_;
  assign new_n_n2015_ = new_n_n543_ | new_n_n1658_;
  assign new_n_n2007_ = new_n_n1178_ | new_n_n509_;
  assign new_n_n1161_ = new_n_n716_ & new_n_n1719_;
  assign new_n_n1988_ = new_n_n1156_ | new_n_n536_;
  assign new_n_n1152_ = new_n_n541_ & new_n_n351_;
  assign new_n_n1147_ = new_n_n545_ & new_n_n514_;
  assign new_n_n1142_ = new_n_n550_ & new_n_n1730_;
  assign new_n_n1108_ = new_n_n83_ & new_n_n583_;
  assign new_n_n1103_ = new_n_n559_ & new_n_n1720_;
  assign new_n_n956_ = new_n_n831_ & new_n_n756_;
  assign new_n_n1776_ = new_n_n845_ | new_n_n1726_;
  assign new_n_n905_ = new_n_n808_ & new_n_n805_;
  assign new_n_n1715_ = ~new_nmusel2_;
  assign new_n_n813_ = ~new_n_n1777_;
  assign new_n_n736_ = ~new_n_n1799_;
  assign new_n_n39_ = ~new_n_n2438_;
  assign new_n_n30_ = ~new_n_n2449_;
  assign new_n_n21_ = ~new_n_n2462_;
  assign new_n_n12_ = ~new_n_n2470_;
  assign new_n_n1585_ = new_n_n26_ & new_n_n840_;
  assign new_n_n2445_ = new_n_n1582_ | new_n_n32_;
  assign new_n_n1451_ = new_n_n219_ & new_n_n1607_;
  assign new_n_n1406_ = new_n_n104_ & new_n_n263_;
  assign new_n_n1400_ = new_n_n267_ & new_n_n268_;
  assign new_n_n1395_ = new_n_n815_ & new_n_n1612_;
  assign new_n_n2203_ = new_n_n1612_ | new_n_n1716_;
  assign new_n_n1364_ = new_n_n304_ & new_n_n305_;
  assign new_n_n1360_ = new_n_n2159_ & new_nb9_;
  assign new_n_n1354_ = new_n_n1714_ & new_n_n315_;
  assign new_n_n2162_ = new_n_n323_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n1344_ = new_n_n1657_ & new_n_n1658_;
  assign new_n_n2151_ = new_n_n1337_ | new_n_n1338_;
  assign new_n_n1332_ = new_n_n1640_ & new_n_n341_;
  assign new_n_n1326_ = new_n_n343_ & new_n_n344_;
  assign new_n_n1305_ = new_n_n369_ & new_n_n351_;
  assign new_n_n2116_ = new_n_n379_ | new_n_n378_;
  assign new_no14_ = new_n_n1295_ | new_n_n388_;
  assign new_n_n2107_ = new_n_n1720_ | new_n_n1630_;
  assign new_n_n1285_ = new_n_n397_ & new_n_n1635_;
  assign new_n_n1279_ = new_n_n405_ & new_n_n1724_;
  assign new_n_n1273_ = new_n_n411_ & new_n_n1628_;
  assign new_n_n2069_ = new_n_n444_ & new_n_n815_;
  assign new_n_n1229_ = new_n_n449_ & new_n_n1719_;
  assign new_n_n1224_ = new_n_n831_ & new_n_n424_;
  assign new_n_n1217_ = new_n_n461_ & new_n_n1646_;
  assign new_n_n2045_ = new_n_n601_ & new_n_n1727_;
  assign new_n_n2002_ = new_n_n523_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n1997_ = new_n_n1719_ | new_n_n1654_;
  assign new_n_n1120_ = new_n_n569_ & new_n_n570_;
  assign new_no8_ = new_n_n1112_ | new_n_n1113_;
  assign new_n_n950_ = new_n_n836_ & new_n_n761_;
  assign new_n_n898_ = new_n_n351_ & new_n_n809_;
  assign new_n_n893_ = new_n_n79_ & new_n_n1714_;
  assign new_n_n888_ = new_n_n824_ & new_n_n1719_;
  assign new_n_n881_ = new_n_n831_ & new_n_n832_;
  assign new_n_n1720_ = ~new_nsh1_;
  assign new_n_n827_ = ~new_n_n1758_;
  assign new_n_n745_ = ~new_n_n1697_;
  assign new_n_n68_ = ~new_n_n2403_;
  assign new_n_n57_ = ~new_n_n2414_;
  assign new_n_n46_ = ~new_n_n2431_;
  assign new_n_n35_ = ~new_n_n2443_;
  assign new_n_n24_ = ~new_n_n2457_;
  assign new_n_n13_ = ~new_n_n2471_;
  assign new_n_n2453_ = new_n_n1609_ | new_n_n1715_;
  assign new_n_n2446_ = new_n_n1714_ | new_n_n815_ | new_n_n258_;
  assign new_n_n2261_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n217_;
  assign new_n_n2219_ = new_n_n1402_ | new_n_n1404_ | new_n_n1403_ | new_n_n1405_;
  assign new_n_n1401_ = new_n_n267_ & new_n_n266_;
  assign new_n_n1394_ = new_n_n282_ & new_n_n1715_;
  assign new_n_n1390_ = new_n_n278_ & new_n_n279_;
  assign new_n_n2178_ = new_n_n1614_ | new_n_n1716_;
  assign new_n_n2173_ = new_n_n1359_ | new_n_n1360_;
  assign new_n_n1353_ = new_n_n1714_ & new_n_n316_;
  assign new_n_n1349_ = new_n_n321_ & new_n_n322_;
  assign new_n_n1343_ = new_n_n1657_ & new_n_n543_;
  assign new_n_n2152_ = new_n_n1658_ & new_n_n543_;
  assign new_n_n2147_ = new_n_n1330_ | new_n_n1331_;
  assign new_n_n2143_ = new_n_n1326_ | new_n_n342_;
  assign new_n_n1304_ = new_n_n369_ & new_n_n370_;
  assign new_n_n2117_ = new_n_n377_ | new_n_n1628_;
  assign new_n_n1295_ = new_n_n389_ & new_n_n1730_;
  assign new_n_n1291_ = new_n_n83_ & new_n_n394_;
  assign new_n_n1284_ = new_n_n397_ & new_n_n398_;
  assign new_n_n1280_ = new_n_n405_ & new_n_n1632_;
  assign new_n_n1267_ = new_n_n416_ & new_n_n1730_;
  assign new_n_n1240_ = new_n_n438_ & new_n_n437_;
  assign new_n_n2063_ = new_n_n1721_ | new_n_n1720_;
  assign new_n_n2058_ = new_n_n1221_ | new_n_n1223_ | new_n_n1222_ | new_n_n1224_;
  assign new_n_n1216_ = new_n_n461_ & new_n_n1724_;
  assign new_n_n1212_ = new_n_n1647_ & new_n_n510_;
  assign new_no10_ = new_n_n1171_ | new_n_n524_;
  assign new_n_n1167_ = new_n_n83_ & new_n_n530_;
  assign new_n_n1119_ = new_n_n1662_ & new_n_n1663_;
  assign new_n_n1114_ = new_n_n574_ & new_n_n575_;
  assign new_n_n1806_ = new_n_n1724_ | new_n_n766_;
  assign new_n_n897_ = new_n_n385_ & new_n_n810_;
  assign new_n_n1764_ = new_n_n890_ | new_n_n892_ | new_n_n891_ | new_n_n893_;
  assign new_n_n1757_ = new_n_n886_ | new_n_n887_;
  assign new_n_n882_ = new_n_n830_ & new_n_n1719_;
  assign new_n_n835_ = ~new_n_n1754_;
  assign new_n_n828_ = ~new_n_n1702_;
  assign new_n_n754_ = ~new_n_n1820_;
  assign new_n_n67_ = ~new_n_n2402_;
  assign new_n_n58_ = ~new_n_n2415_;
  assign new_n_n45_ = ~new_n_n2430_;
  assign new_n_n36_ = ~new_n_n2444_;
  assign new_n_n23_ = ~new_n_n2459_;
  assign new_n_n14_ = ~new_n_n2469_;
  assign new_n_n2460_ = new_n_n1587_ | new_n_n20_;
  assign new_n_n1443_ = new_n_n104_ & new_n_n224_;
  assign new_n_n1405_ = new_n_n1688_ & new_n_n1684_;
  assign new_n_n1399_ = new_n_n269_ & new_n_n1678_;
  assign new_n_n1396_ = new_n_n1670_ & new_n_n598_;
  assign new_n_n2204_ = new_n_n1390_ | new_n_n819_;
  assign new_n_n2177_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n306_;
  assign new_n_n2172_ = new_n_n1355_ | new_n_n1357_ | new_n_n1356_ | new_n_n1358_;
  assign new_n_n2169_ = new_n_n1715_ | new_n_n820_ | new_n_n552_;
  assign new_n_n1350_ = new_n_n321_ & new_n_n1714_;
  assign new_n_n1342_ = new_n_n563_ & new_n_n1658_;
  assign new_n_n1337_ = new_n_n331_ & new_n_n332_;
  assign new_n_n2149_ = new_n_n337_ | new_n_n336_;
  assign new_n_n1327_ = new_n_n341_ & new_n_n376_;
  assign new_n_n2134_ = new_n_n1312_ | new_n_n1311_ | new_n_n1313_ | new_n_n1314_;
  assign new_n_n2128_ = new_n_n1309_ | new_n_n364_;
  assign new_n_n2112_ = new_n_n1721_ | new_n_n1719_;
  assign new_n_n2105_ = new_n_n1290_ | new_n_n395_;
  assign new_n_n1287_ = new_n_n396_ & new_n_n1635_;
  assign new_n_n1281_ = new_n_n853_ & new_n_n1632_;
  assign new_n_n2090_ = new_n_n376_ | new_n_n1640_;
  assign new_no13_ = new_n_n1267_ | new_n_n415_;
  assign new_n_n1239_ = new_n_n438_ & new_n_n1724_;
  assign new_n_n1234_ = new_n_n79_ & new_n_n446_;
  assign new_n_n1225_ = new_n_n451_ & new_n_n1721_;
  assign new_n_n2051_ = new_n_n1216_ | new_n_n913_ | new_n_n1217_ | new_n_n1218_;
  assign new_n_n1213_ = new_n_n466_ & new_n_n467_;
  assign new_n_n1173_ = new_n_n351_ & new_n_n521_;
  assign new_n_n1998_ = new_n_n1167_ | new_n_n529_;
  assign new_n_n940_ = new_n_n730_ & new_n_n731_;
  assign new_n_n1768_ = new_n_n811_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n891_ = new_n_n817_ & new_n_n1714_;
  assign new_n_n1759_ = new_n_n1719_ | new_n_n1718_;
  assign new_n_n1754_ = new_n_n881_ | new_n_n882_;
  assign new_n_n848_ = ~new_n_n1729_;
  assign new_n_n841_ = ~new_n_n1751_;
  assign new_n_n763_ = ~new_n_n1809_;
  assign new_n_n88_ = ~new_n_n2384_;
  assign new_n_n77_ = ~new_n_n2441_;
  assign new_n_n44_ = ~new_n_n2432_;
  assign new_n_n33_ = ~new_n_n2447_;
  assign new_n_n26_ = ~new_n_n2456_;
  assign new_n_n15_ = ~new_n_n2467_;
  assign new_n_n2461_ = new_n_n840_ | new_n_n21_;
  assign new_n_n1438_ = new_n_n1714_ & new_n_n227_;
  assign new_n_n1404_ = new_n_n1688_ & new_n_n675_;
  assign new_n_n2214_ = new_n_n1398_ | new_n_n1399_;
  assign new_n_n2209_ = new_n_n1393_ | new_n_n1395_ | new_n_n1394_ | new_n_n1358_;
  assign new_n_n1391_ = new_n_n1714_ & new_n_n277_;
  assign new_n_n2176_ = new_n_n307_ & new_n_n815_;
  assign new_n_n1359_ = new_n_n104_ & new_n_n313_;
  assign new_n_n2168_ = new_n_n1353_ | new_n_n1354_;
  assign new_n_n1351_ = new_n_n79_ & new_n_n322_;
  assign new_n_n1341_ = new_n_n563_ & new_n_n543_;
  assign new_n_n1338_ = new_n_n1618_ & new_n_n511_;
  assign new_n_n2148_ = new_n_n1332_ | new_n_n376_;
  assign new_n_n1328_ = new_n_n341_ & new_n_n1640_;
  assign new_n_n1314_ = new_n_n833_ & new_n_n836_;
  assign new_n_n2129_ = new_n_n365_ | new_n_n366_;
  assign new_n_n2111_ = new_n_n390_ & new_n_n815_;
  assign new_n_n2106_ = new_n_n1720_ | new_n_n401_;
  assign new_n_n1286_ = new_n_n396_ & new_n_n398_;
  assign new_n_n2097_ = new_n_n1279_ | new_n_n913_ | new_n_n1280_ | new_n_n1281_;
  assign new_n_n2089_ = new_n_n1272_ | new_n_n1273_;
  assign new_n_n2087_ = new_n_n414_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n2072_ = new_n_n1724_ | new_n_n438_;
  assign new_n_n2068_ = new_n_n1232_ | new_n_n1234_ | new_n_n1233_ | new_n_n893_;
  assign new_n_n1230_ = new_n_n449_ & new_n_n1649_;
  assign new_n_n1218_ = new_n_n853_ & new_n_n1646_;
  assign new_n_n2046_ = new_n_n1213_ | new_n_n465_;
  assign new_n_n1172_ = new_n_n385_ & new_n_n522_;
  assign new_n_n1999_ = new_n_n1653_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_ne2_ = new_n_n933_ | new_n_n934_;
  assign new_no1_ = new_n_n896_ | new_n_n812_;
  assign new_n_n892_ = new_n_n79_ & new_n_n818_;
  assign new_n_n1758_ = new_n_n888_ | new_n_n823_;
  assign new_n_n1755_ = new_n_n984_ | new_n_n924_;
  assign new_n_n847_ = ~new_n_n1746_;
  assign new_n_n1724_ = ~new_nopsel2_;
  assign new_n_n1706_ = ~new_n_n2310_;
  assign new_n_n87_ = ~new_n_n2383_;
  assign new_n_n78_ = ~new_n_n1598_;
  assign new_n_n43_ = ~new_n_n2434_;
  assign new_n_n34_ = ~new_n_n2445_;
  assign new_n_n25_ = ~new_n_n2455_;
  assign new_n_n16_ = ~new_n_n2468_;
  assign new_n_n2246_ = new_n_n234_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2199_ = new_n_n284_ & new_n_n1716_ & new_n_n820_;
  assign new_n_n2194_ = new_n_n1715_ | new_n_n820_ | new_n_n488_;
  assign new_n_n1377_ = new_n_n295_ & new_n_n1714_;
  assign new_n_n2175_ = new_n_n1361_ | new_n_n1363_ | new_n_n1362_ | new_n_n893_;
  assign new_n_n1357_ = new_n_n815_ & new_n_n1615_;
  assign new_n_n2166_ = new_n_n1615_ | new_n_n1716_;
  assign new_n_n1347_ = new_n_n848_ & new_n_n1724_;
  assign new_n_n2158_ = new_n_n1345_ | new_n_n1346_;
  assign new_n_n2153_ = new_n_n1339_ | new_n_n1340_;
  assign new_n_n1334_ = new_n_n467_ & new_n_n334_;
  assign new_n_n2144_ = new_n_n1327_ | new_n_n1328_;
  assign new_n_n1320_ = new_n_n385_ & new_n_n352_;
  assign new_n_n1315_ = new_n_n83_ & new_n_n360_;
  assign new_n_n1313_ = new_n_n1721_ & new_n_n836_;
  assign new_n_n2127_ = new_n_n1306_ | new_n_n913_ | new_n_n1307_ | new_n_n1308_;
  assign new_n_n2121_ = new_n_n429_ | new_n_n1638_;
  assign new_ne14_ = new_n_n1298_ | new_n_n1299_;
  assign new_n_n2103_ = new_n_n1720_ & new_n_n1719_;
  assign new_n_n1282_ = new_n_n403_ & new_n_n404_;
  assign new_n_n1275_ = new_n_n1732_ & new_n_n1633_;
  assign new_n_n1268_ = new_n_n385_ & new_n_n413_;
  assign new_n_n1261_ = new_n_n1635_ & new_n_n422_;
  assign new_n_n1253_ = new_n_n425_ & new_n_n426_;
  assign new_n_n1246_ = new_n_n433_ & new_n_n437_;
  assign new_n_n2052_ = new_n_n1219_ | new_n_n458_;
  assign new_n_n2047_ = new_n_n466_ | new_n_n467_;
  assign new_n_n1168_ = new_n_n527_ & new_n_n528_;
  assign new_n_n1793_ = new_n_n927_ | new_n_n929_ | new_n_n928_ | new_n_n893_;
  assign new_n_n876_ = new_n_n836_ & new_n_n837_;
  assign new_n_n1747_ = new_n_n868_ | new_n_n869_;
  assign new_n_n863_ = new_n_n351_ & new_n_n850_;
  assign new_n_n1736_ = new_n_n1735_ & new_n_n860_;
  assign new_n_n860_ = ~new_n_n1658_;
  assign new_n_n855_ = ~new_n_n1747_;
  assign new_n_n779_ = ~new_n_n1804_;
  assign new_n_n89_ = ~new_n_n2381_;
  assign new_n_n86_ = ~new_n_n2390_;
  assign new_n_n75_ = ~new_n_n2393_;
  assign new_n_n64_ = ~new_n_n2407_;
  assign new_n_n53_ = ~new_n_n2422_;
  assign new_n_n28_ = ~new_n_n2453_;
  assign new_n_n17_ = ~new_n_n2464_;
  assign new_n_n2243_ = new_n_n1425_ | new_n_n1427_ | new_n_n1426_ | new_n_n1358_;
  assign new_nb11_ = new_n_n285_ & new_n_n286_;
  assign new_n_n2195_ = new_n_n815_ | new_n_n1713_ | new_n_n1648_;
  assign new_n_n1376_ = new_n_n295_ & new_n_n296_;
  assign new_n_n1363_ = new_n_n79_ & new_n_n309_;
  assign new_n_n1358_ = new_n_n815_ & new_n_n1715_;
  assign new_n_n2165_ = new_n_n1713_ & new_n_n1715_ & new_n_n1714_ & new_n_n319_;
  assign new_n_n1348_ = new_n_n1729_ & new_n_n1730_;
  assign new_n_n1346_ = new_n_n2159_ & new_nb8_;
  assign new_n_n2154_ = new_n_n564_ | new_n_n1617_;
  assign new_n_n1333_ = new_n_n467_ & new_n_n335_;
  assign new_n_n1329_ = new_n_n339_ & new_n_n340_;
  assign new_n_n2139_ = new_n_n353_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n2135_ = new_n_n1315_ | new_n_n359_;
  assign new_n_n1312_ = new_n_n1721_ & new_n_n1719_;
  assign new_n_n1309_ = new_n_n365_ & new_n_n366_;
  assign new_n_n2120_ = new_n_n372_ | new_n_n342_;
  assign new_n_n1300_ = new_n_n383_ & new_n_n380_;
  assign new_n_n2102_ = new_n_n1284_ | new_n_n1286_ | new_n_n1285_ | new_n_n1287_;
  assign new_n_n2098_ = new_n_n1282_ | new_n_n402_;
  assign new_n_n1274_ = new_n_n409_ & new_n_n857_;
  assign new_n_n1269_ = new_n_n351_ & new_n_n412_;
  assign new_n_n2086_ = new_n_n417_ & new_n_n815_;
  assign new_n_n2078_ = new_n_n1251_ | new_n_n1252_;
  assign new_n_n2075_ = new_n_n999_ | new_n_n1245_ | new_n_n1244_ | new_n_n1246_;
  assign new_n_n1219_ = new_n_n459_ & new_n_n460_;
  assign new_n_n1214_ = new_n_n463_ & new_n_n464_;
  assign new_n_n2003_ = new_n_n1172_ | new_n_n1173_;
  assign new_n_n1788_ = new_n_n923_ | new_n_n924_;
  assign new_n_n875_ = new_n_n838_ & new_n_n1721_;
  assign new_n_n1748_ = new_n_n842_ & new_n_n351_;
  assign new_n_n862_ = new_n_n385_ & new_n_n851_;
  assign new_n_n1737_ = new_n_n1688_ & new_n_n2220_;
  assign new_n_n1735_ = ~new_n_n2173_;
  assign new_n_n1730_ = ~new_nopsel3_;
  assign new_n_n788_ = ~new_n_n1654_;
  assign new_n_n1598_ = ~new_nind15_;
  assign new_n_n85_ = ~new_n_n2385_;
  assign new_n_n76_ = ~new_n_n2394_;
  assign new_n_n63_ = ~new_n_n2409_;
  assign new_n_n54_ = ~new_n_n2420_;
  assign new_n_n27_ = ~new_n_n2452_;
  assign new_n_n18_ = ~new_n_n2465_;
  assign new_n_n2238_ = new_n_n1422_ | new_n_n819_;
  assign new_n_n2198_ = new_n_n1385_ | new_n_n1386_;
  assign new_n_n1381_ = new_n_n1714_ & new_n_n289_;
  assign new_n_n2188_ = new_n_n1376_ | new_n_n1378_ | new_n_n1377_ | new_n_n893_;
  assign new_n_n1370_ = new_n_n510_ & new_n_n466_;
  assign new_n_n1362_ = new_n_n308_ & new_n_n1714_;
  assign new_n_n1355_ = new_n_n321_ & new_n_n1615_;
  assign new_n_n2167_ = new_n_n1352_ | new_n_n819_;
  assign new_n_n2161_ = new_n_n1347_ | new_n_n1348_;
  assign new_n_n1345_ = new_n_n104_ & new_n_n327_;
  assign new_n_n1339_ = new_n_n330_ & new_n_n543_;
  assign new_n_n1336_ = new_n_n1620_ & new_n_n334_;
  assign new_n_n2145_ = new_n_n1329_ | new_n_n345_;
  assign new_n_n2140_ = new_n_n1320_ | new_n_n1321_;
  assign new_n_n2136_ = new_n_n1622_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n2133_ = new_n_n1311_ | new_n_n361_;
  assign new_n_n1307_ = new_n_n367_ & new_n_n1625_;
  assign new_n_n2123_ = new_n_n409_ | new_n_n1633_;
  assign new_n_n1301_ = new_n_n383_ & new_n_n342_;
  assign new_n_n1296_ = new_n_n385_ & new_n_n386_;
  assign new_n_n2108_ = new_n_n1291_ | new_n_n393_;
  assign new_n_n1276_ = new_n_n1640_ & new_n_n371_;
  assign new_n_n2088_ = new_n_n1268_ | new_n_n1269_;
  assign new_n_n2085_ = new_n_n1264_ | new_n_n1266_ | new_n_n1265_ | new_n_n893_;
  assign new_n_n1259_ = new_n_n424_ & new_n_n422_;
  assign new_n_n1247_ = new_n_n1640_ & new_n_n432_;
  assign new_n_n2054_ = new_n_n569_ | new_n_n538_ | new_n_n1663_ | new_n_n501_;
  assign new_n_n1215_ = new_n_n463_ & new_n_n351_;
  assign new_n_n918_ = new_n_n790_ & new_n_n789_;
  assign new_n_n1751_ = new_n_n873_ | new_n_n874_;
  assign new_n_n868_ = new_n_n843_ & new_n_n844_;
  assign new_n_n864_ = new_n_n846_ & new_n_n847_;
  assign new_n_n1738_ = new_n_n1734_ & new_n_n859_;
  assign new_n_n90_ = ~new_ninb15_;
  assign new_n_n84_ = ~new_n_n2388_;
  assign new_n_n73_ = ~new_n_n2397_;
  assign new_n_n66_ = ~new_n_n2406_;
  assign new_n_n55_ = ~new_n_n2418_;
  assign new_n_n48_ = ~new_n_n2428_;
  assign new_n_n37_ = ~new_n_n2439_;
  assign new_n_n1386_ = new_n_n2159_ & new_nb11_;
  assign new_n_n2193_ = new_n_n1380_ | new_n_n1381_;
  assign new_n_n1378_ = new_n_n79_ & new_n_n296_;
  assign new_n_n1365_ = new_n_n1714_ & new_n_n303_;
  assign new_n_n1361_ = new_n_n308_ & new_n_n309_;
  assign new_n_n1356_ = new_n_n321_ & new_n_n1715_;
  assign new_n_n1352_ = new_n_n317_ & new_n_n318_;
  assign new_nb8_ = new_n_n324_ & new_n_n325_;
  assign new_n_n2157_ = new_n_n1341_ | new_n_n1343_ | new_n_n1342_ | new_n_n1344_;
  assign new_n_n1340_ = new_n_n330_ & new_n_n1658_;
  assign new_n_n1335_ = new_n_n1620_ & new_n_n335_;
  assign new_n_n2146_ = new_n_n374_ | new_n_n1627_;
  assign new_n_n1321_ = new_n_n351_ & new_n_n586_;
  assign new_n_n1316_ = new_n_n357_ & new_n_n358_;
  assign new_n_n1311_ = new_n_n833_ & new_n_n1719_;
  assign new_n_n1308_ = new_n_n853_ & new_n_n1625_;
  assign new_n_n2122_ = new_n_n2343_ | new_n_n1732_;
  assign new_n_n2115_ = new_n_n1300_ | new_n_n1301_;
  assign new_n_n2113_ = new_n_n387_ | new_n_n853_ | new_n_n1730_;
  assign new_n_n2109_ = new_n_n1629_ | new_n_n820_ | new_n_n1716_ | new_n_n81_;
  assign new_n_n2091_ = new_n_n1274_ | new_n_n1275_;
  assign new_n_n1270_ = new_n_n410_ & new_n_n411_;
  assign new_n_n1266_ = new_n_n79_ & new_n_n419_;
  assign new_n_n1260_ = new_n_n424_ & new_n_n1636_;
  assign new_n_n1254_ = new_n_n425_ & new_n_n836_;
  assign new_n_n2053_ = new_n_n459_ | new_n_n460_;
  assign new_n_n2048_ = new_n_n1214_ | new_n_n1215_;
  assign new_n_n913_ = new_n_n853_ & new_n_n1724_;
  assign new_n_n874_ = new_n_n839_ & new_n_n840_;
  assign new_n_n869_ = new_n_n843_ & new_n_n351_;
  assign new_n_n1744_ = new_n_n862_ | new_n_n863_;
  assign new_n_n1739_ = new_n_n1733_ & new_n_n858_;
  assign new_n_n91_ = ~new_n_n2379_;
  assign new_n_n83_ = ~new_n_n1763_;
  assign new_n_n74_ = ~new_n_n2395_;
  assign new_n_n65_ = ~new_n_n2405_;
  assign new_n_n56_ = ~new_n_n2419_;
  assign new_n_n47_ = ~new_n_n2427_;
  assign new_n_n38_ = ~new_n_n2440_;
endmodule


