// Benchmark "top" written by ABC on Sat Apr  1 09:25:41 2023

module top ( 
    pv28_20_, pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv120_16_, pv120_29_,
    pv168_9_, pv180_10_, pv28_10_, pv56_13_, pv56_22_, pv88_7_, pv88_29_,
    pv120_15_, pv180_4_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_,
    pv120_18_, pv180_5_, pv180_12_, pv192_0_, pv56_15_, pv56_24_, pv88_9_,
    pv88_18_, pv88_27_, pv120_17_, pv168_8_, pv180_6_, pv88_2_, pv88_15_,
    pv88_26_, pv120_12_, pv88_3_, pv88_16_, pv88_25_, pv120_11_, pv180_0_,
    pv56_10_, pv56_21_, pv88_4_, pv88_13_, pv88_24_, pv120_14_, pv126_5_,
    pv180_1_, pv56_11_, pv56_20_, pv88_5_, pv88_14_, pv88_23_, pv120_13_,
    pv180_2_, pv28_8_, pv56_5_, pv88_11_, pv88_22_, pv120_5_, pv132_0_,
    pv156_6_, pv168_1_, pv189_0_, pv28_9_, pv56_4_, pv88_12_, pv88_21_,
    pv120_6_, pv156_5_, pv156_10_, pv168_2_, pv189_1_, pv28_6_, pv56_7_,
    pv88_20_, pv120_3_, pv120_10_, pv156_8_, pv189_2_, pv28_7_, pv56_6_,
    pv88_10_, pv120_4_, pv168_0_, pv28_4_, pv56_9_, pv120_1_, pv168_5_,
    pv28_5_, pv56_8_, pv120_2_, pv156_9_, pv156_14_, pv168_6_, pv28_2_,
    pv156_13_, pv28_3_, pv120_0_, pv156_12_, pv168_4_, pv28_0_, pv186_1_,
    pv28_1_, pv144_4_, pv186_2_, pv144_5_, pv156_0_, pv132_5_, pv144_6_,
    pv56_1_, pv120_9_, pv120_30_, pv132_4_, pv156_2_, pv56_0_, pv88_30_,
    pv132_3_, pv144_8_, pv156_1_, pv28_19_, pv56_3_, pv88_31_, pv120_7_,
    pv132_2_, pv144_9_, pv156_4_, pv56_2_, pv120_8_, pv120_20_, pv132_1_,
    pv186_0_, pv28_17_, pv120_21_, pv126_3_, pv144_10_, pv168_12_,
    pv183_2_, pv28_18_, pv28_27_, pv120_22_, pv126_4_, pv28_15_, pv28_26_,
    pv88_0_, pv120_23_, pv126_1_, pv144_12_, pv168_14_, pv28_16_, pv28_25_,
    pv88_1_, pv120_24_, pv120_31_, pv126_2_, pv168_13_, pv28_13_, pv28_24_,
    pv56_16_, pv56_27_, pv120_25_, pv144_14_, pv180_14_, pv192_2_,
    pv28_14_, pv28_23_, pv56_17_, pv56_26_, pv120_19_, pv120_26_, pv126_0_,
    pv144_0_, pv144_13_, pv180_8_, pv180_13_, pv192_1_, pv28_11_, pv28_22_,
    pv56_18_, pv120_27_, pv144_1_, pv168_10_, pv180_9_, pv183_0_, pv28_12_,
    pv28_21_, pv56_19_, pv120_28_, pv144_2_, pv183_1_,
    pv198_3_, pv198_0_, pv198_2_, pv198_1_, pv194_0_, pv194_1_  );
  input  pv28_20_, pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv120_16_,
    pv120_29_, pv168_9_, pv180_10_, pv28_10_, pv56_13_, pv56_22_, pv88_7_,
    pv88_29_, pv120_15_, pv180_4_, pv56_14_, pv56_25_, pv88_8_, pv88_17_,
    pv88_28_, pv120_18_, pv180_5_, pv180_12_, pv192_0_, pv56_15_, pv56_24_,
    pv88_9_, pv88_18_, pv88_27_, pv120_17_, pv168_8_, pv180_6_, pv88_2_,
    pv88_15_, pv88_26_, pv120_12_, pv88_3_, pv88_16_, pv88_25_, pv120_11_,
    pv180_0_, pv56_10_, pv56_21_, pv88_4_, pv88_13_, pv88_24_, pv120_14_,
    pv126_5_, pv180_1_, pv56_11_, pv56_20_, pv88_5_, pv88_14_, pv88_23_,
    pv120_13_, pv180_2_, pv28_8_, pv56_5_, pv88_11_, pv88_22_, pv120_5_,
    pv132_0_, pv156_6_, pv168_1_, pv189_0_, pv28_9_, pv56_4_, pv88_12_,
    pv88_21_, pv120_6_, pv156_5_, pv156_10_, pv168_2_, pv189_1_, pv28_6_,
    pv56_7_, pv88_20_, pv120_3_, pv120_10_, pv156_8_, pv189_2_, pv28_7_,
    pv56_6_, pv88_10_, pv120_4_, pv168_0_, pv28_4_, pv56_9_, pv120_1_,
    pv168_5_, pv28_5_, pv56_8_, pv120_2_, pv156_9_, pv156_14_, pv168_6_,
    pv28_2_, pv156_13_, pv28_3_, pv120_0_, pv156_12_, pv168_4_, pv28_0_,
    pv186_1_, pv28_1_, pv144_4_, pv186_2_, pv144_5_, pv156_0_, pv132_5_,
    pv144_6_, pv56_1_, pv120_9_, pv120_30_, pv132_4_, pv156_2_, pv56_0_,
    pv88_30_, pv132_3_, pv144_8_, pv156_1_, pv28_19_, pv56_3_, pv88_31_,
    pv120_7_, pv132_2_, pv144_9_, pv156_4_, pv56_2_, pv120_8_, pv120_20_,
    pv132_1_, pv186_0_, pv28_17_, pv120_21_, pv126_3_, pv144_10_,
    pv168_12_, pv183_2_, pv28_18_, pv28_27_, pv120_22_, pv126_4_, pv28_15_,
    pv28_26_, pv88_0_, pv120_23_, pv126_1_, pv144_12_, pv168_14_, pv28_16_,
    pv28_25_, pv88_1_, pv120_24_, pv120_31_, pv126_2_, pv168_13_, pv28_13_,
    pv28_24_, pv56_16_, pv56_27_, pv120_25_, pv144_14_, pv180_14_,
    pv192_2_, pv28_14_, pv28_23_, pv56_17_, pv56_26_, pv120_19_, pv120_26_,
    pv126_0_, pv144_0_, pv144_13_, pv180_8_, pv180_13_, pv192_1_, pv28_11_,
    pv28_22_, pv56_18_, pv120_27_, pv144_1_, pv168_10_, pv180_9_, pv183_0_,
    pv28_12_, pv28_21_, pv56_19_, pv120_28_, pv144_2_, pv183_1_;
  output pv198_3_, pv198_0_, pv198_2_, pv198_1_, pv194_0_, pv194_1_;
  wire new_n_n134_, new_n_n153_, new_n_n128_, new_n_n190_, new_n_n75_,
    new_n_n81_, new_n_n50_, new_n_n82_, new_n_n43_, new_n_n202_,
    new_n_n149_, new_n_n197_, new_n_n102_, new_n_n51_, new_n_n83_,
    new_n_n58_, new_n_n201_, new_n_n122_, new_n_n98_, new_n_n78_,
    new_n_n53_, new_n_n185_, new_n_n55_, new_n_n40_, new_n_n22_,
    new_n_n146_, new_n_n126_, new_n_n96_, new_n_n184_, new_n_n57_,
    new_n_n77_, new_n_n85_, new_n_n52_, new_n_n192_, new_n_n84_,
    new_n_n180_, new_n_n90_, new_n_n111_, new_n_n80_, new_n_n60_,
    new_n_n92_, new_n_n67_, new_n_n203_, new_n_n131_, new_n_n107_,
    new_n_n87_, new_n_n62_, new_n_n187_, new_n_n33_, new_n_n64_,
    new_n_n155_, new_n_n135_, new_n_n105_, new_n_n186_, new_n_n66_,
    new_n_n86_, new_n_n61_, new_n_n161_, new_n_n167_, new_n_n93_,
    new_n_n182_, new_n_n104_, new_n_n45_, new_n_n124_, new_n_n100_,
    new_n_n25_, new_n_n159_, new_n_n171_, new_n_n89_, new_n_n69_,
    new_n_n191_, new_n_n127_, new_n_n115_, new_n_n97_, new_n_n24_,
    new_n_n204_, new_n_n164_, new_n_n71_, new_n_n110_, new_n_n189_,
    new_n_n121_, new_n_n23_, new_n_n165_, new_n_n205_, new_n_n188_,
    new_n_n108_, new_n_n103_, new_n_n170_, new_n_n158_, new_n_n113_,
    new_n_n91_, new_n_n168_, new_n_n162_, new_n_n193_, new_n_n118_,
    new_n_n106_, new_n_n88_, new_n_n206_, new_n_n109_, new_n_n174_,
    new_n_n117_, new_n_n112_, new_n_n94_, new_n_n210_, new_n_n27_,
    new_n_n208_, new_n_n166_, new_n_n26_, new_n_n163_, new_n_n139_,
    new_n_n32_, new_n_n160_, new_n_n209_, new_n_n95_, new_n_n179_,
    new_n_n36_, new_n_n133_, new_n_n211_, new_n_n178_, new_n_n38_,
    new_n_n157_, new_n_n136_, new_n_n138_, new_n_n173_, new_n_n48_,
    new_n_n101_, new_n_n177_, new_n_n154_, new_n_n130_, new_n_n207_,
    new_n_n99_, new_n_n72_, new_n_n41_, new_n_n28_, new_n_n141_,
    new_n_n68_, new_n_n39_, new_n_n151_, new_n_n76_, new_n_n29_,
    new_n_n198_, new_n_n120_, new_n_n183_, new_n_n35_, new_n_n147_,
    new_n_n194_, new_n_n116_, new_n_n65_, new_n_n42_, new_n_n148_,
    new_n_n70_, new_n_n143_, new_n_n123_, new_n_n114_, new_n_n63_,
    new_n_n47_, new_n_n176_, new_n_n73_, new_n_n150_, new_n_n125_,
    new_n_n144_, new_n_n119_, new_n_n59_, new_n_n142_, new_n_n34_,
    new_n_n20_, new_n_n200_, new_n_n129_, new_n_n140_, new_n_n195_,
    new_n_n74_, new_n_n181_, new_n_n44_, new_n_n175_, new_n_n145_,
    new_n_n49_, new_n_n37_, new_n_n21_, new_n_n156_, new_n_n196_,
    new_n_n199_, new_n_n56_, new_n_n172_, new_n_n79_, new_n_n46_,
    new_n_n31_, new_n_n152_, new_n_n132_, new_n_n137_, new_n_n54_,
    new_n_n169_, new_n_n30_, new_nv281_, new_nv285_, new_nv284_,
    new_nv283_, new_nv282_, new_n_n17_, new_n_n18_, new_n_n19_, new_nv286_,
    new_nv207_, new_nv218_, new_n_n11_, new_nv240_, new_nv208_, new_nv217_,
    new_nv230_, new_nv239_, new_nv209_, new_nv220_, new_n_n13_, new_nv238_,
    new_nv210_, new_nv219_, new_n_n12_, new_nv237_, new_n_n16_, new_nv247_,
    new_n_n6_, new_nv269_, new_nv280_, new_nv248_, new_n_n7_, new_nv270_,
    new_nv279_, new_nv249_, new_nv260_, new_nv267_, new_nv278_, new_nv250_,
    new_n_n5_, new_nv268_, new_nv277_, new_nv221_, new_nv232_, new_n_n9_,
    new_nv254_, new_nv265_, new_nv276_, new_nv222_, new_nv231_, new_n_n8_,
    new_nv253_, new_nv266_, new_nv275_, new_nv201_, new_nv212_, new_nv245_,
    new_nv256_, new_nv263_, new_n_n2_, new_nv202_, new_nv211_, new_nv246_,
    new_nv255_, new_nv264_, new_n_n3_, new_nv200_, new_nv203_, new_nv214_,
    new_nv225_, new_nv236_, new_nv261_, new_n_n4_, new_nv199_, new_nv204_,
    new_nv213_, new_nv226_, new_nv235_, new_nv262_, new_nv271_, new_n_n14_,
    new_nv205_, new_nv216_, new_nv223_, new_nv234_, new_nv241_, new_nv252_,
    new_n_n15_, new_nv206_, new_nv215_, new_nv224_, new_nv233_, new_n_n10_,
    new_nv251_;
  assign new_n_n134_ = pv28_20_;
  assign new_n_n153_ = pv56_12_;
  assign new_n_n128_ = pv56_23_;
  assign new_n_n190_ = pv88_6_;
  assign new_n_n75_ = pv88_19_;
  assign new_n_n81_ = pv120_16_;
  assign new_n_n50_ = pv120_29_;
  assign new_n_n82_ = pv168_9_;
  assign new_n_n43_ = pv180_10_;
  assign new_n_n202_ = pv28_10_;
  assign new_n_n149_ = pv56_13_;
  assign new_n_n197_ = pv56_22_;
  assign new_n_n102_ = pv88_7_;
  assign new_n_n51_ = pv88_29_;
  assign new_n_n83_ = pv120_15_;
  assign new_n_n58_ = pv180_4_;
  assign new_n_n201_ = pv56_14_;
  assign new_n_n122_ = pv56_25_;
  assign new_n_n98_ = pv88_8_;
  assign new_n_n78_ = pv88_17_;
  assign new_n_n53_ = pv88_28_;
  assign new_n_n185_ = pv120_18_;
  assign new_n_n55_ = pv180_5_;
  assign new_n_n40_ = pv180_12_;
  assign new_n_n22_ = pv192_0_;
  assign new_n_n146_ = pv56_15_;
  assign new_n_n126_ = pv56_24_;
  assign new_n_n96_ = pv88_9_;
  assign new_n_n184_ = pv88_18_;
  assign new_n_n57_ = pv88_27_;
  assign new_n_n77_ = pv120_17_;
  assign new_n_n85_ = pv168_8_;
  assign new_n_n52_ = pv180_6_;
  assign new_n_n192_ = pv88_2_;
  assign new_n_n84_ = pv88_15_;
  assign new_n_n180_ = pv88_26_;
  assign new_n_n90_ = pv120_12_;
  assign new_n_n111_ = pv88_3_;
  assign new_n_n80_ = pv88_16_;
  assign new_n_n60_ = pv88_25_;
  assign new_n_n92_ = pv120_11_;
  assign new_n_n67_ = pv180_0_;
  assign new_n_n203_ = pv56_10_;
  assign new_n_n131_ = pv56_21_;
  assign new_n_n107_ = pv88_4_;
  assign new_n_n87_ = pv88_13_;
  assign new_n_n62_ = pv88_24_;
  assign new_n_n187_ = pv120_14_;
  assign new_n_n33_ = pv126_5_;
  assign new_n_n64_ = pv180_1_;
  assign new_n_n155_ = pv56_11_;
  assign new_n_n135_ = pv56_20_;
  assign new_n_n105_ = pv88_5_;
  assign new_n_n186_ = pv88_14_;
  assign new_n_n66_ = pv88_23_;
  assign new_n_n86_ = pv120_13_;
  assign new_n_n61_ = pv180_2_;
  assign new_n_n161_ = pv28_8_;
  assign new_n_n167_ = pv56_5_;
  assign new_n_n93_ = pv88_11_;
  assign new_n_n182_ = pv88_22_;
  assign new_n_n104_ = pv120_5_;
  assign new_n_n45_ = pv132_0_;
  assign new_n_n124_ = pv156_6_;
  assign new_n_n100_ = pv168_1_;
  assign new_n_n25_ = pv189_0_;
  assign new_n_n159_ = pv28_9_;
  assign new_n_n171_ = pv56_4_;
  assign new_n_n89_ = pv88_12_;
  assign new_n_n69_ = pv88_21_;
  assign new_n_n191_ = pv120_6_;
  assign new_n_n127_ = pv156_5_;
  assign new_n_n115_ = pv156_10_;
  assign new_n_n97_ = pv168_2_;
  assign new_n_n24_ = pv189_1_;
  assign pv198_3_ = new_n_n16_;
  assign new_n_n204_ = pv28_6_;
  assign new_n_n164_ = pv56_7_;
  assign new_n_n71_ = pv88_20_;
  assign new_n_n110_ = pv120_3_;
  assign new_n_n189_ = pv120_10_;
  assign new_n_n121_ = pv156_8_;
  assign new_n_n23_ = pv189_2_;
  assign new_n_n165_ = pv28_7_;
  assign new_n_n205_ = pv56_6_;
  assign new_n_n188_ = pv88_10_;
  assign new_n_n108_ = pv120_4_;
  assign new_n_n103_ = pv168_0_;
  assign new_n_n170_ = pv28_4_;
  assign new_n_n158_ = pv56_9_;
  assign new_n_n113_ = pv120_1_;
  assign new_n_n91_ = pv168_5_;
  assign pv198_0_ = new_n_n19_;
  assign new_n_n168_ = pv28_5_;
  assign new_n_n162_ = pv56_8_;
  assign new_n_n193_ = pv120_2_;
  assign new_n_n118_ = pv156_9_;
  assign new_n_n106_ = pv156_14_;
  assign new_n_n88_ = pv168_6_;
  assign new_n_n206_ = pv28_2_;
  assign new_n_n109_ = pv156_13_;
  assign pv198_2_ = new_n_n17_;
  assign new_n_n174_ = pv28_3_;
  assign new_n_n117_ = pv120_0_;
  assign new_n_n112_ = pv156_12_;
  assign new_n_n94_ = pv168_4_;
  assign pv198_1_ = new_n_n18_;
  assign new_n_n210_ = pv28_0_;
  assign new_n_n27_ = pv186_1_;
  assign new_n_n208_ = pv28_1_;
  assign new_n_n166_ = pv144_4_;
  assign new_n_n26_ = pv186_2_;
  assign new_n_n163_ = pv144_5_;
  assign new_n_n139_ = pv156_0_;
  assign new_n_n32_ = pv132_5_;
  assign new_n_n160_ = pv144_6_;
  assign new_n_n209_ = pv56_1_;
  assign new_n_n95_ = pv120_9_;
  assign new_n_n179_ = pv120_30_;
  assign new_n_n36_ = pv132_4_;
  assign new_n_n133_ = pv156_2_;
  assign new_n_n211_ = pv56_0_;
  assign new_n_n178_ = pv88_30_;
  assign new_n_n38_ = pv132_3_;
  assign new_n_n157_ = pv144_8_;
  assign new_n_n136_ = pv156_1_;
  assign new_n_n138_ = pv28_19_;
  assign new_n_n173_ = pv56_3_;
  assign new_n_n48_ = pv88_31_;
  assign new_n_n101_ = pv120_7_;
  assign new_n_n177_ = pv132_2_;
  assign new_n_n154_ = pv144_9_;
  assign new_n_n130_ = pv156_4_;
  assign new_n_n207_ = pv56_2_;
  assign new_n_n99_ = pv120_8_;
  assign new_n_n72_ = pv120_20_;
  assign new_n_n41_ = pv132_1_;
  assign new_n_n28_ = pv186_0_;
  assign new_n_n141_ = pv28_17_;
  assign new_n_n68_ = pv120_21_;
  assign new_n_n39_ = pv126_3_;
  assign new_n_n151_ = pv144_10_;
  assign new_n_n76_ = pv168_12_;
  assign new_n_n29_ = pv183_2_;
  assign pv194_0_ = new_n_n15_;
  assign new_n_n198_ = pv28_18_;
  assign new_n_n120_ = pv28_27_;
  assign new_n_n183_ = pv120_22_;
  assign new_n_n35_ = pv126_4_;
  assign new_n_n147_ = pv28_15_;
  assign new_n_n194_ = pv28_26_;
  assign new_n_n116_ = pv88_0_;
  assign new_n_n65_ = pv120_23_;
  assign new_n_n42_ = pv126_1_;
  assign new_n_n148_ = pv144_12_;
  assign new_n_n70_ = pv168_14_;
  assign new_n_n143_ = pv28_16_;
  assign new_n_n123_ = pv28_25_;
  assign new_n_n114_ = pv88_1_;
  assign new_n_n63_ = pv120_24_;
  assign new_n_n47_ = pv120_31_;
  assign new_n_n176_ = pv126_2_;
  assign new_n_n73_ = pv168_13_;
  assign pv194_1_ = new_n_n14_;
  assign new_n_n150_ = pv28_13_;
  assign new_n_n125_ = pv28_24_;
  assign new_n_n144_ = pv56_16_;
  assign new_n_n119_ = pv56_27_;
  assign new_n_n59_ = pv120_25_;
  assign new_n_n142_ = pv144_14_;
  assign new_n_n34_ = pv180_14_;
  assign new_n_n20_ = pv192_2_;
  assign new_n_n200_ = pv28_14_;
  assign new_n_n129_ = pv28_23_;
  assign new_n_n140_ = pv56_17_;
  assign new_n_n195_ = pv56_26_;
  assign new_n_n74_ = pv120_19_;
  assign new_n_n181_ = pv120_26_;
  assign new_n_n44_ = pv126_0_;
  assign new_n_n175_ = pv144_0_;
  assign new_n_n145_ = pv144_13_;
  assign new_n_n49_ = pv180_8_;
  assign new_n_n37_ = pv180_13_;
  assign new_n_n21_ = pv192_1_;
  assign new_n_n156_ = pv28_11_;
  assign new_n_n196_ = pv28_22_;
  assign new_n_n199_ = pv56_18_;
  assign new_n_n56_ = pv120_27_;
  assign new_n_n172_ = pv144_1_;
  assign new_n_n79_ = pv168_10_;
  assign new_n_n46_ = pv180_9_;
  assign new_n_n31_ = pv183_0_;
  assign new_n_n152_ = pv28_12_;
  assign new_n_n132_ = pv28_21_;
  assign new_n_n137_ = pv56_19_;
  assign new_n_n54_ = pv120_28_;
  assign new_n_n169_ = pv144_2_;
  assign new_n_n30_ = pv183_1_;
  assign new_nv281_ = new_n_n7_ & new_n_n25_;
  assign new_nv285_ = new_n_n21_ & new_n_n3_ & new_n_n22_;
  assign new_nv284_ = new_n_n4_ & new_n_n22_;
  assign new_nv283_ = new_n_n23_ & new_n_n5_ & new_n_n24_ & new_n_n25_;
  assign new_nv282_ = new_n_n24_ & new_n_n6_ & new_n_n25_;
  assign new_n_n17_ = new_nv283_ | new_nv282_ | new_nv281_ | new_nv247_ | new_nv245_ | new_nv207_ | new_nv246_;
  assign new_n_n18_ = new_nv280_ | new_nv279_ | new_nv278_ | new_nv232_ | new_nv230_ | new_nv203_ | new_nv231_;
  assign new_n_n19_ = new_nv277_ | new_nv276_ | new_nv275_ | new_nv217_ | new_nv215_ | new_nv199_ | new_nv216_;
  assign new_nv286_ = new_n_n20_ & new_n_n2_ & new_n_n21_ & new_n_n22_;
  assign new_nv207_ = new_n_n190_ & new_n_n191_;
  assign new_nv218_ = new_n_n166_ & new_n_n165_ & new_n_n164_;
  assign new_n_n11_ = new_nv224_ | new_nv225_ | new_nv226_ | new_nv202_;
  assign new_nv240_ = new_n_n109_ & new_n_n107_ & new_n_n112_ & new_n_n108_;
  assign new_nv208_ = new_n_n188_ & new_n_n189_;
  assign new_nv217_ = new_n_n169_ & new_n_n168_ & new_n_n175_ & new_n_n167_ & new_n_n172_;
  assign new_nv230_ = new_n_n139_ & new_n_n138_ & new_n_n137_;
  assign new_nv239_ = new_n_n112_ & new_n_n111_ & new_n_n110_;
  assign new_nv209_ = new_n_n186_ & new_n_n187_;
  assign new_nv220_ = new_n_n160_ & new_n_n159_ & new_n_n166_ & new_n_n158_ & new_n_n163_;
  assign new_n_n13_ = new_nv218_ | new_nv219_ | new_nv220_ | new_nv200_;
  assign new_nv238_ = new_n_n115_ & new_n_n114_ & new_n_n121_ & new_n_n113_ & new_n_n118_;
  assign new_nv210_ = new_n_n184_ & new_n_n185_;
  assign new_nv219_ = new_n_n163_ & new_n_n161_ & new_n_n166_ & new_n_n162_;
  assign new_n_n12_ = new_nv221_ | new_nv222_ | new_nv223_ | new_nv201_;
  assign new_nv237_ = new_n_n118_ & new_n_n116_ & new_n_n121_ & new_n_n117_;
  assign new_n_n16_ = new_nv286_ | new_nv285_ | new_nv284_ | new_nv262_ | new_nv260_ | new_nv211_ | new_nv261_;
  assign new_nv247_ = new_n_n97_ & new_n_n96_ & new_n_n103_ & new_n_n95_ & new_n_n100_;
  assign new_n_n6_ = new_nv251_ | new_nv252_ | new_nv253_ | new_nv209_;
  assign new_nv269_ = new_n_n40_ & new_n_n39_ & new_n_n38_;
  assign new_nv280_ = new_n_n26_ & new_n_n8_ & new_n_n27_ & new_n_n28_;
  assign new_nv248_ = new_n_n94_ & new_n_n93_ & new_n_n92_;
  assign new_n_n7_ = new_nv248_ | new_nv249_ | new_nv250_ | new_nv208_;
  assign new_nv270_ = new_n_n37_ & new_n_n35_ & new_n_n40_ & new_n_n36_;
  assign new_nv279_ = new_n_n27_ & new_n_n9_ & new_n_n28_;
  assign new_nv249_ = new_n_n91_ & new_n_n89_ & new_n_n94_ & new_n_n90_;
  assign new_nv260_ = new_n_n67_ & new_n_n66_ & new_n_n65_;
  assign new_nv267_ = new_n_n46_ & new_n_n44_ & new_n_n49_ & new_n_n45_;
  assign new_nv278_ = new_n_n10_ & new_n_n28_;
  assign new_nv250_ = new_n_n88_ & new_n_n87_ & new_n_n94_ & new_n_n86_ & new_n_n91_;
  assign new_n_n5_ = new_nv254_ | new_nv255_ | new_nv256_ | new_nv210_;
  assign new_nv268_ = new_n_n43_ & new_n_n42_ & new_n_n49_ & new_n_n41_ & new_n_n46_;
  assign new_nv277_ = new_n_n29_ & new_n_n11_ & new_n_n30_ & new_n_n31_;
  assign new_nv221_ = new_n_n157_ & new_n_n156_ & new_n_n155_;
  assign new_nv232_ = new_n_n133_ & new_n_n132_ & new_n_n139_ & new_n_n131_ & new_n_n136_;
  assign new_n_n9_ = new_nv236_ | new_nv237_ | new_nv238_ | new_nv205_;
  assign new_nv254_ = new_n_n76_ & new_n_n75_ & new_n_n74_;
  assign new_nv265_ = new_n_n52_ & new_n_n51_ & new_n_n58_ & new_n_n50_ & new_n_n55_;
  assign new_nv276_ = new_n_n30_ & new_n_n12_ & new_n_n31_;
  assign new_nv222_ = new_n_n154_ & new_n_n152_ & new_n_n157_ & new_n_n153_;
  assign new_nv231_ = new_n_n136_ & new_n_n134_ & new_n_n139_ & new_n_n135_;
  assign new_n_n8_ = new_nv239_ | new_nv240_ | new_nv241_ | new_nv206_;
  assign new_nv253_ = new_n_n79_ & new_n_n78_ & new_n_n85_ & new_n_n77_ & new_n_n82_;
  assign new_nv266_ = new_n_n49_ & new_n_n48_ & new_n_n47_;
  assign new_nv275_ = new_n_n13_ & new_n_n31_;
  assign new_nv201_ = new_n_n202_ & new_n_n203_;
  assign new_nv212_ = new_n_n180_ & new_n_n181_;
  assign new_nv245_ = new_n_n103_ & new_n_n102_ & new_n_n101_;
  assign new_nv256_ = new_n_n70_ & new_n_n69_ & new_n_n76_ & new_n_n68_ & new_n_n73_;
  assign new_nv263_ = new_n_n58_ & new_n_n57_ & new_n_n56_;
  assign new_n_n2_ = new_nv269_ | new_nv270_ | new_nv271_ | new_nv214_;
  assign new_nv202_ = new_n_n200_ & new_n_n201_;
  assign new_nv211_ = new_n_n182_ & new_n_n183_;
  assign new_nv246_ = new_n_n100_ & new_n_n98_ & new_n_n103_ & new_n_n99_;
  assign new_nv255_ = new_n_n73_ & new_n_n71_ & new_n_n76_ & new_n_n72_;
  assign new_nv264_ = new_n_n55_ & new_n_n53_ & new_n_n58_ & new_n_n54_;
  assign new_n_n3_ = new_nv266_ | new_nv267_ | new_nv268_ | new_nv213_;
  assign new_nv200_ = new_n_n204_ & new_n_n205_;
  assign new_nv203_ = new_n_n198_ & new_n_n199_;
  assign new_nv214_ = new_n_n176_ & new_n_n177_;
  assign new_nv225_ = new_n_n145_ & new_n_n143_ & new_n_n148_ & new_n_n144_;
  assign new_nv236_ = new_n_n121_ & new_n_n120_ & new_n_n119_;
  assign new_nv261_ = new_n_n64_ & new_n_n62_ & new_n_n67_ & new_n_n63_;
  assign new_n_n4_ = new_nv263_ | new_nv264_ | new_nv265_ | new_nv212_;
  assign new_nv199_ = new_n_n206_ & new_n_n207_;
  assign new_nv204_ = new_n_n196_ & new_n_n197_;
  assign new_nv213_ = new_n_n178_ & new_n_n179_;
  assign new_nv226_ = new_n_n142_ & new_n_n141_ & new_n_n148_ & new_n_n140_ & new_n_n145_;
  assign new_nv235_ = new_n_n124_ & new_n_n123_ & new_n_n130_ & new_n_n122_ & new_n_n127_;
  assign new_nv262_ = new_n_n61_ & new_n_n60_ & new_n_n67_ & new_n_n59_ & new_n_n64_;
  assign new_nv271_ = new_n_n34_ & new_n_n33_ & new_n_n40_ & new_n_n32_ & new_n_n37_;
  assign new_n_n14_ = new_n_n208_ & new_n_n209_;
  assign new_nv205_ = new_n_n194_ & new_n_n195_;
  assign new_nv216_ = new_n_n172_ & new_n_n170_ & new_n_n175_ & new_n_n171_;
  assign new_nv223_ = new_n_n151_ & new_n_n150_ & new_n_n157_ & new_n_n149_ & new_n_n154_;
  assign new_nv234_ = new_n_n127_ & new_n_n125_ & new_n_n130_ & new_n_n126_;
  assign new_nv241_ = new_n_n106_ & new_n_n105_ & new_n_n112_ & new_n_n104_ & new_n_n109_;
  assign new_nv252_ = new_n_n82_ & new_n_n80_ & new_n_n85_ & new_n_n81_;
  assign new_n_n15_ = new_n_n210_ & new_n_n211_;
  assign new_nv206_ = new_n_n192_ & new_n_n193_;
  assign new_nv215_ = new_n_n175_ & new_n_n174_ & new_n_n173_;
  assign new_nv224_ = new_n_n148_ & new_n_n147_ & new_n_n146_;
  assign new_nv233_ = new_n_n130_ & new_n_n129_ & new_n_n128_;
  assign new_n_n10_ = new_nv233_ | new_nv234_ | new_nv235_ | new_nv204_;
  assign new_nv251_ = new_n_n85_ & new_n_n84_ & new_n_n83_;
endmodule


