// Benchmark "top" written by ABC on Fri Mar 31 12:11:33 2023

module top ( 
    pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1, pf4, pr,
    pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0, pf3,
    pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, pk3, px, ph1, pi0, pj3, pk2, py, ph2, pi3, pj0, pk1, pz, ph3,
    pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pl1, pm0, pn3, po2, pl2, pm3,
    pn0, po1, pl3, pm2, pn1, po0, pq1, pr2, ps3, pp1, pr3, ps2, pb, pp2,
    pq3, pr0, ps1, pc, pp3, pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1,
    pu0, pv3, pw2, pf, pt2, pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0,
    py1, pz2, pi, px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl,
    pm, pn, po,
    pe5, pf6, pg7, pd5, pf7, pg6, pd6, pe7, pg5, pd7, pe6, pf5, pa5, pb6,
    pc7, pb7, pc6, pa7, pc5, pa6, pb5, pl4, pm5, pn6, po7, pa8, pl5, pm4,
    pn7, po6, pb8, pl6, pm7, pn4, po5, pc8, pl7, pm6, pn5, po4, pi5, pj6,
    pk7, ph5, pi4, pj7, pk6, ph6, pi7, pj4, pk5, ph7, pi6, pj5, pk4, pt4,
    pu5, pv6, pw7, pt5, pu4, pv7, pw6, pt6, pu7, pv4, pw5, pt7, pu6, pv5,
    pw4, pp4, pq5, pr6, ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7,
    pq6, pr5, ps4, px4, py5, pz6, px5, py4, pz7, px6, py7, pz4, px7, py6,
    pz5  );
  input  pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1,
    pf4, pr, pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0,
    pf3, pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw,
    ph0, pi1, pj2, pk3, px, ph1, pi0, pj3, pk2, py, ph2, pi3, pj0, pk1, pz,
    ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pl1, pm0, pn3, po2, pl2,
    pm3, pn0, po1, pl3, pm2, pn1, po0, pq1, pr2, ps3, pp1, pr3, ps2, pb,
    pp2, pq3, pr0, ps1, pc, pp3, pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe,
    pt1, pu0, pv3, pw2, pf, pt2, pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph,
    px0, py1, pz2, pi, px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1,
    pl, pm, pn, po;
  output pe5, pf6, pg7, pd5, pf7, pg6, pd6, pe7, pg5, pd7, pe6, pf5, pa5, pb6,
    pc7, pb7, pc6, pa7, pc5, pa6, pb5, pl4, pm5, pn6, po7, pa8, pl5, pm4,
    pn7, po6, pb8, pl6, pm7, pn4, po5, pc8, pl7, pm6, pn5, po4, pi5, pj6,
    pk7, ph5, pi4, pj7, pk6, ph6, pi7, pj4, pk5, ph7, pi6, pj5, pk4, pt4,
    pu5, pv6, pw7, pt5, pu4, pv7, pw6, pt6, pu7, pv4, pw5, pt7, pu6, pv5,
    pw4, pp4, pq5, pr6, ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7,
    pq6, pr5, ps4, px4, py5, pz6, px5, py4, pz7, px6, py7, pz4, px7, py6,
    pz5;
  wire new_na1_, new_nb2_, new_nc3_, new_nd4_, new_np_, new_na0_, new_nb3_,
    new_nc2_, new_ne4_, new_nq_, new_na3_, new_nb0_, new_nc1_, new_nf4_,
    new_nr_, new_na2_, new_nb1_, new_nc0_, new_ng4_, new_ns_, new_nd0_,
    new_ne1_, new_nf2_, new_ng3_, new_nt_, new_na4_, new_nd1_, new_ne0_,
    new_nf3_, new_ng2_, new_nu_, new_nb4_, new_nd2_, new_ne3_, new_nf0_,
    new_ng1_, new_nv_, new_nc4_, new_nd3_, new_ne2_, new_nf1_, new_ng0_,
    new_nw_, new_nh0_, new_ni1_, new_nj2_, new_nk3_, new_nx_, new_nh1_,
    new_ni0_, new_nj3_, new_nk2_, new_ny_, new_nh2_, new_ni3_, new_nj0_,
    new_nk1_, new_nz_, new_nh3_, new_ni2_, new_nj1_, new_nk0_, new_nh4_,
    new_nl0_, new_nm1_, new_nn2_, new_no3_, new_nl1_, new_nm0_, new_nn3_,
    new_no2_, new_nl2_, new_nm3_, new_nn0_, new_no1_, new_nl3_, new_nm2_,
    new_nn1_, new_no0_, new_nq1_, new_nr2_, new_ns3_, new_np1_, new_nr3_,
    new_ns2_, new_nb_, new_np2_, new_nq3_, new_nr0_, new_ns1_, new_nc_,
    new_np3_, new_nq2_, new_nr1_, new_ns0_, new_nd_, new_nt0_, new_nu1_,
    new_nv2_, new_nw3_, new_ne_, new_nt1_, new_nu0_, new_nv3_, new_nw2_,
    new_nf_, new_nt2_, new_nu3_, new_nv0_, new_nw1_, new_ng_, new_nt3_,
    new_nu2_, new_nv1_, new_nw0_, new_nh_, new_nx0_, new_ny1_, new_nz2_,
    new_ni_, new_nx1_, new_ny0_, new_nz3_, new_nj_, new_nx2_, new_ny3_,
    new_nz0_, new_nk_, new_nx3_, new_ny2_, new_nz1_, new_nl_, new_nm_,
    new_nn_, new_no_, new_nl4_, new_nu4_, new_nf5_, new_nq5_, new_n_n928_,
    new_nh6_, new_n_n898_, new_n_n889_, new_n_n880_, new_n_n872_, new_nt6_,
    new_n_n857_, new_n_n850_, new_n_n842_, new_n_n811_, new_nr7_,
    new_n_n795_, new_nx7_, new_n_n777_, new_n_n768_, new_n_n760_,
    new_n_n752_, new_n_n747_, new_nq12_, new_n_n730_, new_n_n722_,
    new_n_n687_, new_n_n678_, new_n_n669_, new_nq14_, new_n_n652_,
    new_n_n643_, new_n_n634_, new_n_n608_, new_n_n599_, new_n_n590_,
    new_n_n583_, new_n_n573_, new_n_n569_, new_n_n561_, new_ny16_,
    new_ng18_, new_nq18_, new_n_n543_, new_ne19_, new_nu19_, new_na20_,
    new_n_n523_, new_n_n516_, new_ny20_, new_n_n501_, new_n_n494_,
    new_n_n488_, new_n_n481_, new_n_n474_, new_n_n467_, new_n_n460_,
    new_n_n453_, new_n_n446_, new_n_n439_, new_n_n432_, new_n_n425_,
    new_n_n418_, new_n_n411_, new_n_n404_, new_n_n397_, new_n_n390_,
    new_nq24_, new_na25_, new_n_n371_, new_n_n365_, new_n_n356_,
    new_n_n345_, new_n_n334_, new_n_n323_, new_n_n312_, new_n_n301_,
    new_n_n268_, new_n_n257_, new_n_n246_, new_n_n235_, new_n_n224_,
    new_n_n213_, new_n_n202_, new_n_n158_, new_n_n147_, new_n_n136_,
    new_n_n125_, new_n_n114_, new_n_n103_, new_n_n935_, new_nv4_, new_ne5_,
    new_nr5_, new_n_n929_, new_n_n914_, new_nj6_, new_n_n890_, new_n_n879_,
    new_np6_, new_n_n864_, new_n_n858_, new_n_n849_, new_n_n843_,
    new_n_n810_, new_n_n803_, new_nv7_, new_n_n787_, new_n_n776_, new_na8_,
    new_n_n759_, new_n_n753_, new_n_n746_, new_n_n739_, new_n_n729_,
    new_n_n723_, new_n_n686_, new_n_n679_, new_nm14_, new_n_n661_,
    new_n_n651_, new_n_n644_, new_n_n626_, new_n_n607_, new_n_n600_,
    new_n_n589_, new_n_n584_, new_n_n572_, new_np16_, new_n_n560_,
    new_n_n555_, new_n_n553_, new_np18_, new_n_n542_, new_nc19_,
    new_n_n536_, new_n_n531_, new_nj20_, new_np20_, new_n_n502_, new_ng21_,
    new_n_n495_, new_n_n487_, new_nt21_, new_n_n473_, new_nd22_,
    new_n_n459_, new_nn22_, new_n_n445_, new_nx22_, new_n_n438_,
    new_n_n424_, new_nm23_, new_n_n410_, new_nw23_, new_n_n396_,
    new_n_n391_, new_nr24_, new_nz24_, new_n_n370_, new_nm25_, new_n_n355_,
    new_n_n346_, new_n_n333_, new_n_n324_, new_n_n311_, new_n_n302_,
    new_n_n278_, new_n_n256_, new_n_n247_, new_n_n234_, new_n_n225_,
    new_n_n212_, new_n_n203_, new_n_n157_, new_n_n148_, new_n_n135_,
    new_n_n126_, new_n_n113_, new_n_n104_, new_n_n933_, new_ns4_, new_nd5_,
    new_n_n921_, new_n_n915_, new_n_n897_, new_n_n887_, new_n_n882_,
    new_n_n873_, new_n_n863_, new_n_n856_, new_n_n851_, new_n_n844_,
    new_n_n826_, new_nm7_, new_n_n794_, new_n_n785_, new_n_n779_,
    new_n_n769_, new_n_n762_, new_n_n754_, new_n_n745_, new_n_n737_,
    new_n_n732_, new_nb13_, new_nc14_, new_n_n680_, new_n_n668_,
    new_n_n659_, new_n_n653_, new_na15_, new_n_n618_, new_n_n609_,
    new_nw15_, new_nc16_, new_n_n581_, new_n_n575_, new_n_n570_, new_nr17_,
    new_n_n554_, new_no18_, new_nx18_, new_n_n537_, new_nr19_, new_ny19_,
    new_n_n522_, new_n_n510_, new_ne21_, new_np21_, new_nu21_, new_n_n475_,
    new_n_n468_, new_nj22_, new_no22_, new_n_n447_, new_n_n440_, new_ni23_,
    new_nn23_, new_n_n412_, new_n_n405_, new_nc24_, new_nj24_, new_no24_,
    new_n_n387_, new_nh25_, new_nn25_, new_n_n358_, new_n_n347_,
    new_n_n332_, new_n_n321_, new_n_n314_, new_n_n303_, new_n_n277_,
    new_n_n266_, new_n_n248_, new_n_n233_, new_n_n222_, new_n_n215_,
    new_n_n204_, new_n_n178_, new_n_n167_, new_n_n134_, new_n_n123_,
    new_n_n116_, new_n_n105_, new_n_n934_, new_nt4_, new_nc5_, new_n_n920_,
    new_nd6_, new_n_n896_, new_n_n888_, new_n_n881_, new_n_n874_, new_nu6_,
    new_nx6_, new_na7_, new_nd7_, new_n_n825_, new_n_n818_, new_n_n793_,
    new_n_n786_, new_n_n778_, new_n_n770_, new_n_n761_, new_nz11_,
    new_n_n744_, new_n_n738_, new_n_n731_, new_n_n724_, new_n_n688_,
    new_ng14_, new_n_n667_, new_n_n660_, new_nu14_, new_n_n645_,
    new_n_n610_, new_ns15_, new_n_n601_, new_nd16_, new_n_n582_,
    new_n_n574_, new_no16_, new_nu17_, new_ne18_, new_nf18_, new_n_n541_,
    new_nh19_, new_ns19_, new_n_n532_, new_n_n515_, new_n_n509_,
    new_n_n503_, new_nq21_, new_n_n480_, new_ny21_, new_n_n469_, new_nk22_,
    new_n_n452_, new_ns22_, new_n_n441_, new_nj23_, new_n_n417_, new_nr23_,
    new_n_n406_, new_nd24_, new_nh24_, new_np24_, new_ny24_, new_ni25_,
    new_n_n364_, new_n_n357_, new_n_n348_, new_n_n331_, new_n_n322_,
    new_n_n313_, new_n_n304_, new_n_n276_, new_n_n267_, new_n_n258_,
    new_n_n232_, new_n_n223_, new_n_n214_, new_n_n205_, new_n_n177_,
    new_n_n168_, new_n_n133_, new_n_n124_, new_n_n115_, new_n_n106_,
    new_nn4_, new_nm5_, new_n_n930_, new_n_n922_, new_nc6_, new_n_n895_,
    new_nl6_, new_nn6_, new_n_n869_, new_n_n867_, new_n_n860_, new_nz6_,
    new_n_n845_, new_n_n824_, new_n_n816_, new_n_n808_, new_ns7_, new_ny7_,
    new_n_n771_, new_nc8_, new_nk12_, new_nl12_, new_no12_, new_n_n734_,
    new_n_n725_, new_n_n684_, new_n_n675_, new_nk14_, new_n_n664_,
    new_n_n655_, new_n_n646_, new_nu15_, new_n_n596_, new_n_n593_,
    new_n_n587_, new_n_n577_, new_nn16_, new_n_n551_, new_nr18_,
    new_n_n538_, new_no19_, new_n_n533_, new_nh21_, new_n_n493_,
    new_n_n477_, new_n_n470_, new_n_n437_, new_n_n430_, new_n_n407_,
    new_n_n395_, new_n_n385_, new_n_n376_, new_n_n330_, new_n_n319_,
    new_n_n297_, new_n_n286_, new_n_n231_, new_n_n220_, new_n_n209_,
    new_n_n198_, new_n_n187_, new_n_n132_, new_n_n121_, new_n_n110_,
    new_n_n99_, new_n_n8_, new_nm4_, new_nn5_, new_n_n931_, new_ny5_,
    new_nb6_, new_n_n894_, new_n_n886_, new_n_n876_, new_n_n870_, new_ns6_,
    new_nv6_, new_n_n852_, new_n_n846_, new_nk7_, new_n_n817_, new_n_n807_,
    new_n_n800_, new_n_n780_, new_n_n772_, new_n_n756_, new_nj12_,
    new_nn12_, new_n_n741_, new_n_n733_, new_n_n726_, new_n_n683_,
    new_n_n676_, new_n_n672_, new_no14_, new_n_n654_, new_n_n647_,
    new_n_n604_, new_ny15_, new_na16_, new_n_n588_, new_n_n576_, new_nm16_,
    new_n_n550_, new_n_n547_, new_n_n545_, new_nq19_, new_nx19_, new_ni21_,
    new_nm21_, new_n_n476_, new_nc22_, new_n_n436_, new_ne23_, new_n_n413_,
    new_n_n389_, new_n_n384_, new_n_n377_, new_n_n329_, new_n_n320_,
    new_n_n296_, new_n_n287_, new_n_n230_, new_n_n221_, new_n_n199_,
    new_n_n197_, new_n_n188_, new_n_n131_, new_n_n122_, new_n_n109_,
    new_n_n100_, new_nw4_, new_nh5_, new_no5_, new_nw5_, new_nx5_,
    new_n_n916_, new_n_n893_, new_n_n884_, new_n_n878_, new_nq6_,
    new_n_n866_, new_nw6_, new_n_n854_, new_nc7_, new_n_n823_, new_nn7_,
    new_n_n809_, new_n_n801_, new_nu7_, new_n_n788_, new_n_n758_,
    new_ni12_, new_n_n749_, new_n_n740_, new_nw12_, new_na13_, new_n_n685_,
    new_ni14_, new_n_n671_, new_n_n662_, new_ns14_, new_n_n648_,
    new_n_n606_, new_n_n597_, new_n_n592_, new_n_n585_, new_n_n579_,
    new_nl16_, new_nh18_, new_n_n548_, new_n_n544_, new_nb19_, new_n_n534_,
    new_n_n500_, new_nl21_, new_n_n489_, new_n_n482_, new_ny22_, new_nd23_,
    new_n_n419_, new_ns24_, new_n_n386_, new_n_n378_, new_n_n310_,
    new_n_n299_, new_n_n288_, new_n_n229_, new_n_n211_, new_n_n200_,
    new_n_n130_, new_n_n119_, new_n_n112_, new_n_n101_, new_nx4_, new_ng5_,
    new_np5_, new_nv5_, new_n_n923_, new_n_n917_, new_n_n892_, new_n_n885_,
    new_n_n877_, new_n_n871_, new_n_n865_, new_n_n859_, new_n_n853_,
    new_n_n847_, new_n_n822_, new_n_n815_, new_np7_, new_n_n802_,
    new_n_n796_, new_n_n789_, new_n_n757_, new_nc12_, new_n_n748_,
    new_np12_, new_n_n735_, new_nz12_, new_ne14_, new_n_n677_, new_n_n670_,
    new_n_n663_, new_n_n656_, new_ny14_, new_n_n605_, new_n_n598_,
    new_n_n591_, new_n_n586_, new_n_n578_, new_nj16_, new_n_n552_,
    new_n_n549_, new_nw18_, new_na19_, new_nn19_, new_n_n499_, new_nk21_,
    new_no21_, new_n_n483_, new_nz22_, new_n_n431_, new_nh23_, new_nb25_,
    new_nc25_, new_n_n379_, new_n_n309_, new_n_n300_, new_n_n298_,
    new_n_n219_, new_n_n210_, new_n_n201_, new_n_n129_, new_n_n120_,
    new_n_n111_, new_n_n102_, new_ni5_, new_nt5_, new_n_n925_, new_na6_,
    new_ng6_, new_n_n901_, new_n_n848_, new_n_n838_, new_ni7_, new_n_n720_,
    new_n_n711_, new_n_n702_, new_n_n693_, new_nc15_, new_n_n632_,
    new_n_n623_, new_n_n614_, new_n_n566_, new_n_n559_, new_ne17_,
    new_ny17_, new_nk18_, new_n_n521_, new_n_n514_, new_na21_, new_n_n496_,
    new_n_n490_, new_np22_, new_nu22_, new_n_n434_, new_n_n427_,
    new_n_n420_, new_nt24_, new_nd25_, new_n_n373_, new_nl25_, new_n_n359_,
    new_n_n293_, new_n_n282_, new_n_n271_, new_n_n260_, new_n_n249_,
    new_n_n194_, new_n_n183_, new_n_n172_, new_n_n161_, new_n_n150_,
    new_n_n139_, new_n_n4_, new_nj5_, new_ns5_, new_n_n924_, new_n_n918_,
    new_n_n909_, new_n_n902_, new_ny6_, new_n_n837_, new_n_n830_,
    new_n_n719_, new_n_n712_, new_n_n701_, new_n_n694_, new_n_n640_,
    new_ng15_, new_n_n622_, new_n_n615_, new_n_n565_, new_nt16_, new_ng17_,
    new_nx17_, new_nu18_, new_n_n528_, new_n_n513_, new_n_n507_, new_nj21_,
    new_n_n491_, new_n_n451_, new_nt22_, new_n_n433_, new_n_n428_,
    new_n_n414_, new_nk24_, new_n_n381_, new_n_n374_, new_n_n366_,
    new_n_n360_, new_n_n292_, new_n_n283_, new_n_n270_, new_n_n261_,
    new_n_n239_, new_n_n193_, new_n_n184_, new_n_n171_, new_n_n162_,
    new_n_n149_, new_n_n140_, new_n_n5_, new_nk5_, new_nu5_, new_n_n927_,
    new_n_n919_, new_n_n911_, new_n_n903_, new_n_n861_, new_n_n839_,
    new_n_n831_, new_n_n718_, new_n_n709_, new_n_n704_, new_n_n695_,
    new_n_n682_, new_n_n639_, new_n_n630_, new_nk15_, new_n_n616_,
    new_n_n603_, new_n_n594_, new_nq16_, new_n_n557_, new_nc17_, new_nw17_,
    new_ni18_, new_n_n546_, new_n_n527_, new_n_n520_, new_n_n508_,
    new_n_n498_, new_nn21_, new_n_n464_, new_n_n457_, new_nb23_, new_ng23_,
    new_nv23_, new_n_n394_, new_n_n383_, new_n_n375_, new_n_n350_,
    new_n_n339_, new_n_n295_, new_n_n284_, new_n_n269_, new_n_n251_,
    new_n_n240_, new_n_n196_, new_n_n185_, new_n_n170_, new_n_n159_,
    new_n_n152_, new_n_n141_, new_n_n6_, new_nl5_, new_n_n932_,
    new_n_n926_, new_nz5_, new_n_n910_, new_ni6_, new_n_n868_, new_nf7_,
    new_n_n832_, new_n_n717_, new_n_n710_, new_n_n703_, new_n_n696_,
    new_n_n674_, new_n_n638_, new_n_n631_, new_n_n624_, new_no15_,
    new_n_n602_, new_n_n595_, new_nr16_, new_n_n558_, new_nd17_, new_nv17_,
    new_nj18_, new_ns18_, new_nf20_, new_nl20_, new_ns20_, new_n_n497_,
    new_n_n492_, new_nh22_, new_n_n458_, new_n_n435_, new_n_n429_,
    new_n_n401_, new_na24_, new_n_n382_, new_nf25_, new_n_n349_,
    new_n_n340_, new_n_n294_, new_n_n285_, new_n_n259_, new_n_n250_,
    new_n_n241_, new_n_n195_, new_n_n186_, new_n_n169_, new_n_n160_,
    new_n_n151_, new_n_n142_, new_n_n7_, new_n_n937_, new_nq4_, new_nb5_,
    new_n_n912_, new_n_n904_, new_no6_, new_n_n841_, new_nh7_, new_nm13_,
    new_n_n708_, new_n_n699_, new_n_n690_, new_n_n666_, new_n_n637_,
    new_ni15_, new_n_n620_, new_n_n611_, new_nf16_, new_nh16_, new_n_n564_,
    new_nw16_, new_nj17_, new_nd18_, new_n_n540_, new_nj19_, new_n_n535_,
    new_n_n526_, new_nn20_, new_n_n511_, new_n_n504_, new_n_n486_,
    new_n_n479_, new_n_n472_, new_n_n465_, new_n_n463_, new_n_n456_,
    new_n_n449_, new_n_n442_, new_n_n423_, new_n_n416_, new_n_n409_,
    new_n_n402_, new_n_n400_, new_n_n393_, new_nm24_, new_nx24_, new_nj25_,
    new_n_n363_, new_n_n352_, new_n_n341_, new_n_n338_, new_n_n327_,
    new_n_n316_, new_n_n305_, new_n_n289_, new_n_n275_, new_n_n264_,
    new_n_n253_, new_n_n242_, new_n_n228_, new_n_n217_, new_n_n206_,
    new_n_n190_, new_n_n179_, new_n_n176_, new_n_n165_, new_n_n154_,
    new_n_n143_, new_n_n118_, new_n_n107_, new_n_n0_, new_nj4_, new_nr4_,
    new_na5_, new_nf6_, new_n_n905_, new_nm6_, new_n_n840_, new_n_n833_,
    new_n_n716_, new_ns13_, new_n_n698_, new_n_n691_, new_n_n658_,
    new_ne15_, new_n_n629_, new_n_n619_, new_n_n612_, new_ng16_,
    new_n_n580_, new_ns16_, new_nv16_, new_nk17_, new_nb18_, new_nz18_,
    new_ni19_, new_nd20_, new_n_n525_, new_n_n519_, new_nw20_, new_nc21_,
    new_n_n485_, new_nv21_, new_n_n471_, new_nf22_, new_n_n462_, new_nm22_,
    new_n_n448_, new_nw22_, new_n_n422_, new_no23_, new_n_n408_, new_ny23_,
    new_n_n399_, new_nf24_, new_nn24_, new_nw24_, new_n_n369_, new_no25_,
    new_n_n351_, new_n_n342_, new_n_n337_, new_n_n328_, new_n_n315_,
    new_n_n306_, new_n_n279_, new_n_n274_, new_n_n265_, new_n_n252_,
    new_n_n243_, new_n_n238_, new_n_n216_, new_n_n207_, new_n_n189_,
    new_n_n180_, new_n_n175_, new_n_n166_, new_n_n153_, new_n_n144_,
    new_n_n117_, new_n_n108_, new_n_n1_, new_n_n936_, new_no4_, new_nz4_,
    new_ne6_, new_n_n906_, new_n_n891_, new_n_n715_, new_n_n706_,
    new_nw13_, new_n_n692_, new_n_n650_, new_n_n636_, new_n_n627_,
    new_n_n621_, new_nq15_, new_n_n571_, new_n_n567_, new_n_n563_,
    new_n_n556_, new_nh17_, new_na18_, new_n_n539_, new_nv19_, new_n_n529_,
    new_nh20_, new_n_n517_, new_nu20_, new_n_n505_, new_ns21_, new_nx21_,
    new_nz21_, new_ne22_, new_n_n461_, new_n_n454_, new_n_n450_,
    new_n_n443_, new_nc23_, new_nl23_, new_nq23_, new_ns23_, new_nx23_,
    new_n_n398_, new_ng24_, new_n_n388_, new_nv24_, new_n_n380_,
    new_n_n372_, new_n_n368_, new_n_n361_, new_n_n354_, new_n_n343_,
    new_n_n336_, new_n_n325_, new_n_n318_, new_n_n307_, new_n_n291_,
    new_n_n280_, new_n_n273_, new_n_n262_, new_n_n255_, new_n_n244_,
    new_n_n237_, new_n_n226_, new_n_n208_, new_n_n192_, new_n_n181_,
    new_n_n174_, new_n_n163_, new_n_n156_, new_n_n145_, new_n_n138_,
    new_n_n127_, new_n_n2_, new_nk4_, new_np4_, new_ny4_, new_n_n913_,
    new_n_n907_, new_n_n899_, new_n_n714_, new_n_n707_, new_n_n700_,
    new_na14_, new_n_n642_, new_n_n635_, new_n_n628_, new_nm15_,
    new_n_n613_, new_ni16_, new_n_n568_, new_n_n562_, new_nx16_, new_ni17_,
    new_nz17_, new_nl19_, new_nw19_, new_n_n530_, new_n_n524_, new_n_n518_,
    new_n_n512_, new_n_n506_, new_n_n484_, new_n_n478_, new_na22_,
    new_n_n466_, new_ni22_, new_n_n455_, new_nr22_, new_n_n444_,
    new_n_n426_, new_n_n421_, new_n_n415_, new_nt23_, new_n_n403_,
    new_nb24_, new_n_n392_, new_nl24_, new_nu24_, new_ne25_, new_ng25_,
    new_n_n367_, new_n_n362_, new_n_n353_, new_n_n344_, new_n_n335_,
    new_n_n326_, new_n_n317_, new_n_n308_, new_n_n290_, new_n_n281_,
    new_n_n272_, new_n_n263_, new_n_n254_, new_n_n245_, new_n_n236_,
    new_n_n227_, new_n_n218_, new_n_n191_, new_n_n182_, new_n_n173_,
    new_n_n164_, new_n_n155_, new_n_n146_, new_n_n137_, new_n_n128_,
    new_n_n3_, new_n_n93_, new_n_n82_, new_n_n71_, new_n_n60_, new_n_n49_,
    new_n_n94_, new_n_n81_, new_n_n72_, new_n_n59_, new_n_n50_, new_n_n95_,
    new_n_n80_, new_n_n69_, new_n_n62_, new_n_n51_, new_n_n96_, new_n_n79_,
    new_n_n70_, new_n_n61_, new_n_n52_, new_ni4_, new_n_n835_, new_nj7_,
    new_n_n705_, new_ny13_, new_n_n617_, new_n_n97_, new_n_n42_,
    new_n_n31_, new_n_n20_, new_n_n9_, new_n_n834_, new_n_n827_, new_nu13_,
    new_n_n697_, new_n_n625_, new_n_n98_, new_n_n41_, new_n_n32_,
    new_n_n19_, new_n_n10_, new_n_n908_, new_n_n836_, new_n_n828_,
    new_nc13_, new_nq13_, new_n_n633_, new_n_n40_, new_n_n29_, new_n_n22_,
    new_n_n11_, new_n_n900_, new_ng7_, new_n_n829_, new_n_n721_,
    new_n_n713_, new_n_n641_, new_n_n39_, new_n_n30_, new_n_n21_,
    new_n_n12_, new_nk6_, new_n_n821_, new_n_n813_, new_n_n805_, new_nt7_,
    new_n_n736_, new_n_n727_, new_n_n649_, new_n_n68_, new_n_n57_,
    new_n_n46_, new_n_n35_, new_n_n24_, new_n_n13_, new_n_n883_, new_nl7_,
    new_n_n814_, new_n_n804_, new_n_n797_, new_nr12_, new_n_n728_,
    new_n_n657_, new_n_n67_, new_n_n58_, new_n_n45_, new_n_n36_,
    new_n_n23_, new_n_n14_, new_n_n875_, new_n_n820_, new_no7_,
    new_n_n806_, new_n_n798_, new_n_n751_, new_n_n742_, new_n_n665_,
    new_n_n88_, new_n_n77_, new_n_n44_, new_n_n33_, new_n_n26_, new_n_n15_,
    new_nr6_, new_n_n819_, new_n_n812_, new_nq7_, new_n_n799_, new_n_n750_,
    new_n_n743_, new_n_n673_, new_n_n87_, new_n_n78_, new_n_n43_,
    new_n_n34_, new_n_n25_, new_n_n16_, new_n_n862_, new_nw7_, new_n_n783_,
    new_n_n774_, new_n_n764_, new_n_n763_, new_ny11_, new_n_n681_,
    new_n_n89_, new_n_n86_, new_n_n75_, new_n_n64_, new_n_n53_, new_n_n28_,
    new_n_n17_, new_n_n855_, new_n_n792_, new_n_n784_, new_n_n773_,
    new_n_n765_, new_nb8_, new_n_n755_, new_n_n689_, new_n_n90_,
    new_n_n85_, new_n_n76_, new_n_n63_, new_n_n54_, new_n_n27_, new_n_n18_,
    new_nb7_, new_n_n791_, new_n_n781_, new_n_n775_, new_n_n766_,
    new_n_n91_, new_n_n84_, new_n_n73_, new_n_n66_, new_n_n55_, new_n_n48_,
    new_n_n37_, new_ne7_, new_n_n790_, new_n_n782_, new_nz7_, new_n_n767_,
    new_n_n92_, new_n_n83_, new_n_n74_, new_n_n65_, new_n_n56_, new_n_n47_,
    new_n_n38_;
  assign new_na1_ = pa1;
  assign new_nb2_ = pb2;
  assign new_nc3_ = pc3;
  assign new_nd4_ = pd4;
  assign pe5 = new_ne5_;
  assign pf6 = new_nf6_;
  assign pg7 = new_ng7_;
  assign new_np_ = pp;
  assign new_na0_ = pa0;
  assign new_nb3_ = pb3;
  assign new_nc2_ = pc2;
  assign pd5 = new_nd5_;
  assign new_ne4_ = pe4;
  assign pf7 = new_nf7_;
  assign pg6 = new_ng6_;
  assign new_nq_ = pq;
  assign new_na3_ = pa3;
  assign new_nb0_ = pb0;
  assign new_nc1_ = pc1;
  assign pd6 = new_nd6_;
  assign pe7 = new_ne7_;
  assign new_nf4_ = pf4;
  assign pg5 = new_ng5_;
  assign new_nr_ = pr;
  assign new_na2_ = pa2;
  assign new_nb1_ = pb1;
  assign new_nc0_ = pc0;
  assign pd7 = new_nd7_;
  assign pe6 = new_ne6_;
  assign pf5 = new_nf5_;
  assign new_ng4_ = pg4;
  assign new_ns_ = ps;
  assign pa5 = new_na5_;
  assign pb6 = new_nb6_;
  assign pc7 = new_nc7_;
  assign new_nd0_ = pd0;
  assign new_ne1_ = pe1;
  assign new_nf2_ = pf2;
  assign new_ng3_ = pg3;
  assign new_nt_ = pt;
  assign new_na4_ = pa4;
  assign pb7 = new_nb7_;
  assign pc6 = new_nc6_;
  assign new_nd1_ = pd1;
  assign new_ne0_ = pe0;
  assign new_nf3_ = pf3;
  assign new_ng2_ = pg2;
  assign new_nu_ = pu;
  assign pa7 = new_na7_;
  assign new_nb4_ = pb4;
  assign pc5 = new_nc5_;
  assign new_nd2_ = pd2;
  assign new_ne3_ = pe3;
  assign new_nf0_ = pf0;
  assign new_ng1_ = pg1;
  assign new_nv_ = pv;
  assign pa6 = new_na6_;
  assign pb5 = new_nb5_;
  assign new_nc4_ = pc4;
  assign new_nd3_ = pd3;
  assign new_ne2_ = pe2;
  assign new_nf1_ = pf1;
  assign new_ng0_ = pg0;
  assign new_nw_ = pw;
  assign new_nh0_ = ph0;
  assign new_ni1_ = pi1;
  assign new_nj2_ = pj2;
  assign new_nk3_ = pk3;
  assign pl4 = new_nl4_;
  assign pm5 = new_nm5_;
  assign pn6 = new_nn6_;
  assign po7 = new_no7_;
  assign new_nx_ = px;
  assign pa8 = new_na8_;
  assign new_nh1_ = ph1;
  assign new_ni0_ = pi0;
  assign new_nj3_ = pj3;
  assign new_nk2_ = pk2;
  assign pl5 = new_nl5_;
  assign pm4 = new_nm4_;
  assign pn7 = new_nn7_;
  assign po6 = new_no6_;
  assign new_ny_ = py;
  assign pb8 = new_nb8_;
  assign new_nh2_ = ph2;
  assign new_ni3_ = pi3;
  assign new_nj0_ = pj0;
  assign new_nk1_ = pk1;
  assign pl6 = new_nl6_;
  assign pm7 = new_nm7_;
  assign pn4 = new_nn4_;
  assign po5 = new_no5_;
  assign new_nz_ = pz;
  assign pc8 = new_nc8_;
  assign new_nh3_ = ph3;
  assign new_ni2_ = pi2;
  assign new_nj1_ = pj1;
  assign new_nk0_ = pk0;
  assign pl7 = new_nl7_;
  assign pm6 = new_nm6_;
  assign pn5 = new_nn5_;
  assign po4 = new_no4_;
  assign new_nh4_ = ph4;
  assign pi5 = new_ni5_;
  assign pj6 = new_nj6_;
  assign pk7 = new_nk7_;
  assign new_nl0_ = pl0;
  assign new_nm1_ = pm1;
  assign new_nn2_ = pn2;
  assign new_no3_ = po3;
  assign ph5 = new_nh5_;
  assign pi4 = new_ni4_;
  assign pj7 = new_nj7_;
  assign pk6 = new_nk6_;
  assign new_nl1_ = pl1;
  assign new_nm0_ = pm0;
  assign new_nn3_ = pn3;
  assign new_no2_ = po2;
  assign ph6 = new_nh6_;
  assign pi7 = new_ni7_;
  assign pj4 = new_nj4_;
  assign pk5 = new_nk5_;
  assign new_nl2_ = pl2;
  assign new_nm3_ = pm3;
  assign new_nn0_ = pn0;
  assign new_no1_ = po1;
  assign ph7 = new_nh7_;
  assign pi6 = new_ni6_;
  assign pj5 = new_nj5_;
  assign pk4 = new_nk4_;
  assign new_nl3_ = pl3;
  assign new_nm2_ = pm2;
  assign new_nn1_ = pn1;
  assign new_no0_ = po0;
  assign new_nq1_ = pq1;
  assign new_nr2_ = pr2;
  assign new_ns3_ = ps3;
  assign pt4 = new_nt4_;
  assign pu5 = new_nu5_;
  assign pv6 = new_nv6_;
  assign pw7 = new_nw7_;
  assign new_np1_ = pp1;
  assign new_nr3_ = pr3;
  assign new_ns2_ = ps2;
  assign pt5 = new_nt5_;
  assign pu4 = new_nu4_;
  assign pv7 = new_nv7_;
  assign pw6 = new_nw6_;
  assign new_nb_ = pb;
  assign new_np2_ = pp2;
  assign new_nq3_ = pq3;
  assign new_nr0_ = pr0;
  assign new_ns1_ = ps1;
  assign pt6 = new_nt6_;
  assign pu7 = new_nu7_;
  assign pv4 = new_nv4_;
  assign pw5 = new_nw5_;
  assign new_nc_ = pc;
  assign new_np3_ = pp3;
  assign new_nq2_ = pq2;
  assign new_nr1_ = pr1;
  assign new_ns0_ = ps0;
  assign pt7 = new_nt7_;
  assign pu6 = new_nu6_;
  assign pv5 = new_nv5_;
  assign pw4 = new_nw4_;
  assign new_nd_ = pd;
  assign pp4 = new_np4_;
  assign pq5 = new_nq5_;
  assign pr6 = new_nr6_;
  assign ps7 = new_ns7_;
  assign new_nt0_ = pt0;
  assign new_nu1_ = pu1;
  assign new_nv2_ = pv2;
  assign new_nw3_ = pw3;
  assign new_ne_ = pe;
  assign pp5 = new_np5_;
  assign pq4 = new_nq4_;
  assign pr7 = new_nr7_;
  assign ps6 = new_ns6_;
  assign new_nt1_ = pt1;
  assign new_nu0_ = pu0;
  assign new_nv3_ = pv3;
  assign new_nw2_ = pw2;
  assign new_nf_ = pf;
  assign pp6 = new_np6_;
  assign pq7 = new_nq7_;
  assign pr4 = new_nr4_;
  assign ps5 = new_ns5_;
  assign new_nt2_ = pt2;
  assign new_nu3_ = pu3;
  assign new_nv0_ = pv0;
  assign new_nw1_ = pw1;
  assign new_ng_ = pg;
  assign pp7 = new_np7_;
  assign pq6 = new_nq6_;
  assign pr5 = new_nr5_;
  assign ps4 = new_ns4_;
  assign new_nt3_ = pt3;
  assign new_nu2_ = pu2;
  assign new_nv1_ = pv1;
  assign new_nw0_ = pw0;
  assign new_nh_ = ph;
  assign new_nx0_ = px0;
  assign new_ny1_ = py1;
  assign new_nz2_ = pz2;
  assign new_ni_ = pi;
  assign new_nx1_ = px1;
  assign new_ny0_ = py0;
  assign new_nz3_ = pz3;
  assign new_nj_ = pj;
  assign new_nx2_ = px2;
  assign new_ny3_ = py3;
  assign new_nz0_ = pz0;
  assign new_nk_ = pk;
  assign new_nx3_ = px3;
  assign new_ny2_ = py2;
  assign new_nz1_ = pz1;
  assign new_nl_ = pl;
  assign px4 = new_nx4_;
  assign py5 = new_ny5_;
  assign pz6 = new_nz6_;
  assign new_nm_ = pm;
  assign px5 = new_nx5_;
  assign py4 = new_ny4_;
  assign pz7 = new_nz7_;
  assign new_nn_ = pn;
  assign px6 = new_nx6_;
  assign py7 = new_ny7_;
  assign pz4 = new_nz4_;
  assign new_no_ = po;
  assign px7 = new_nx7_;
  assign py6 = new_ny6_;
  assign pz5 = new_nz5_;
  assign new_nl4_ = new_n_n933_ | new_n_n934_;
  assign new_nu4_ = new_n_n15_ & new_n_n175_;
  assign new_nf5_ = new_n_n26_ & new_n_n175_;
  assign new_nq5_ = new_n_n37_ & new_n_n175_;
  assign new_n_n928_ = new_n_n336_ & new_nb2_ & new_n_n132_;
  assign new_nh6_ = new_n_n904_ | new_n_n906_ | new_n_n905_ | new_n_n907_;
  assign new_n_n898_ = new_n_n71_ & new_n_n67_ & new_n_n175_;
  assign new_n_n889_ = new_n_n71_ & new_np2_ & new_n_n175_;
  assign new_n_n880_ = new_n_n74_ & new_nr2_ & new_n_n175_;
  assign new_n_n872_ = new_n_n77_ & new_nu2_;
  assign new_nt6_ = new_n_n863_ | new_n_n864_;
  assign new_n_n857_ = new_n_n84_ & new_nh_;
  assign new_n_n850_ = new_n_n88_ & new_nf3_;
  assign new_n_n842_ = new_n_n92_ & new_n_n175_ & new_n_n91_;
  assign new_n_n811_ = new_nc_ & new_n_n175_ & new_n_n113_;
  assign new_nr7_ = new_n_n802_ | new_n_n801_ | new_n_n800_;
  assign new_n_n795_ = new_n_n125_ & new_ny3_;
  assign new_nx7_ = new_n_n785_ | new_n_n783_ | new_n_n782_ | new_n_n781_ | new_n_n784_ | new_n_n786_;
  assign new_n_n777_ = new_n_n335_ & new_n_n129_ & new_n_n132_;
  assign new_n_n768_ = new_n_n338_ & new_nf4_ & new_n_n132_;
  assign new_n_n760_ = new_n_n134_ & new_ng4_ & new_n_n132_;
  assign new_n_n752_ = new_n_n136_ & new_n_n137_;
  assign new_n_n747_ = new_n_n325_ & new_n_n141_;
  assign new_nq12_ = new_n_n738_ | new_n_n737_ | new_n_n736_;
  assign new_n_n730_ = new_n_n173_ & new_n_n225_ & new_n_n145_;
  assign new_n_n722_ = new_n_n147_ & new_nr2_;
  assign new_n_n687_ = new_n_n286_ & new_n_n157_;
  assign new_n_n678_ = new_n_n296_ & new_n_n156_;
  assign new_n_n669_ = new_ni_ & new_n_n151_ & new_nr_;
  assign new_nq14_ = new_n_n657_ | new_n_n659_ | new_n_n658_ | new_n_n660_;
  assign new_n_n652_ = new_n_n249_ & new_n_n165_;
  assign new_n_n643_ = new_n_n260_ & new_n_n160_;
  assign new_n_n634_ = new_n_n270_ & new_nb0_;
  assign new_n_n608_ = new_n_n305_ & new_n_n165_;
  assign new_n_n599_ = new_n_n315_ & new_n_n163_;
  assign new_n_n590_ = new_n_n327_ & new_n_n166_;
  assign new_n_n583_ = new_n_n173_ & new_n_n168_ & new_n_n170_;
  assign new_n_n573_ = new_nq12_ & new_n_n318_ & new_n_n172_;
  assign new_n_n569_ = new_n_n225_ & new_n_n325_;
  assign new_n_n561_ = new_nc0_ & new_n_n181_;
  assign new_ny16_ = new_n_n335_ | new_n_n332_ | new_n_n184_;
  assign new_ng18_ = new_n_n553_ | new_ni18_;
  assign new_nq18_ = new_n_n549_ | new_n_n548_ | new_n_n547_;
  assign new_n_n543_ = new_no2_ & new_n_n223_ & new_n_n210_;
  assign new_ne19_ = new_n_n329_ & new_nx1_;
  assign new_nu19_ = new_n_n363_ | new_n_n219_ | new_n_n536_;
  assign new_na20_ = new_ny1_ | new_n_n530_ | new_n_n529_;
  assign new_n_n523_ = new_nf_ & new_n_n235_ & new_n_n231_;
  assign new_n_n516_ = new_n_n234_ & new_n_n244_;
  assign new_ny20_ = new_ny1_ | new_n_n508_ | new_n_n507_;
  assign new_n_n501_ = new_nf_ & new_n_n243_ & new_nh_;
  assign new_n_n494_ = new_nd_ & new_n_n329_ & new_n_n250_;
  assign new_n_n488_ = new_n_n255_ & new_ne_;
  assign new_n_n481_ = new_n_n260_ & new_ne_;
  assign new_n_n474_ = new_n_n265_ & new_ne_;
  assign new_n_n467_ = new_n_n270_ & new_ne_;
  assign new_n_n460_ = new_n_n275_ & new_ne_;
  assign new_n_n453_ = new_n_n280_ & new_ne_;
  assign new_n_n446_ = new_n_n285_ & new_ne_;
  assign new_n_n439_ = new_n_n290_ & new_ne_;
  assign new_n_n432_ = new_n_n295_ & new_ne_;
  assign new_n_n425_ = new_n_n300_ & new_ne_;
  assign new_n_n418_ = new_n_n305_ & new_ne_;
  assign new_n_n411_ = new_n_n310_ & new_ne_;
  assign new_n_n404_ = new_n_n315_ & new_ne_;
  assign new_n_n397_ = new_n_n320_ & new_ne_;
  assign new_n_n390_ = new_nd_ & new_n_n329_ & new_n_n328_;
  assign new_nq24_ = new_ne4_ & new_n_n346_ & new_nc4_;
  assign new_na25_ = new_na4_ & new_nb4_ & new_n_n343_;
  assign new_n_n371_ = new_nl2_ & new_n_n353_;
  assign new_n_n365_ = new_nj2_ & new_nl2_ & new_n_n359_;
  assign new_n_n356_ = ~new_nm25_;
  assign new_n_n345_ = ~new_nc25_;
  assign new_n_n334_ = ~new_ns24_;
  assign new_n_n323_ = ~new_nj2_;
  assign new_n_n312_ = ~new_nw3_;
  assign new_n_n301_ = ~new_nb1_;
  assign new_n_n268_ = ~new_nf22_;
  assign new_n_n257_ = ~new_nl3_;
  assign new_n_n246_ = ~new_nj3_;
  assign new_n_n235_ = ~new_nh_;
  assign new_n_n224_ = ~new_nq2_;
  assign new_n_n213_ = ~new_nn25_;
  assign new_n_n202_ = ~new_nl0_;
  assign new_n_n158_ = ~new_nt_;
  assign new_n_n147_ = ~new_nc13_;
  assign new_n_n136_ = ~new_no0_;
  assign new_n_n125_ = ~new_nj24_;
  assign new_n_n114_ = ~new_nl23_;
  assign new_n_n103_ = ~new_nn22_;
  assign new_n_n935_ = new_n_n325_ & new_n_n6_ & new_nw12_;
  assign new_nv4_ = new_n_n16_ & new_n_n175_;
  assign new_ne5_ = new_n_n25_ & new_n_n175_;
  assign new_nr5_ = new_n_n38_ & new_n_n175_;
  assign new_n_n929_ = new_n_n45_ & new_nb2_ & new_n_n132_;
  assign new_n_n914_ = new_n_n325_ & new_n_n175_ & new_nx19_;
  assign new_nj6_ = new_n_n896_ | new_n_n894_ | new_n_n893_ | new_n_n892_ | new_n_n895_ | new_n_n897_;
  assign new_n_n890_ = new_n_n69_ & new_np2_ & new_n_n175_;
  assign new_n_n879_ = new_nx1_ & new_n_n73_ & new_n_n175_;
  assign new_np6_ = new_n_n871_ | new_n_n872_;
  assign new_n_n864_ = new_n_n81_ & new_ny2_;
  assign new_n_n858_ = new_n_n84_ & new_nb3_;
  assign new_n_n849_ = new_n_n88_ & new_nh_;
  assign new_n_n843_ = new_n_n121_ & new_n_n175_ & new_n_n91_;
  assign new_n_n810_ = new_n_n121_ & new_n_n175_ & new_n_n113_;
  assign new_n_n803_ = new_n_n118_ & new_n_n175_ & new_n_n117_;
  assign new_nv7_ = new_n_n793_ | new_n_n794_;
  assign new_n_n787_ = new_n_n331_ & new_n_n127_ & new_n_n132_;
  assign new_n_n776_ = new_n_n333_ & new_n_n129_ & new_n_n132_;
  assign new_na8_ = new_n_n767_ | new_n_n765_ | new_n_n764_ | new_n_n763_ | new_n_n766_ | new_n_n768_;
  assign new_n_n759_ = new_n_n186_ & new_n_n133_ & new_n_n132_;
  assign new_n_n753_ = new_n_n136_ & new_nx1_;
  assign new_n_n746_ = new_n_n169_ & new_n_n138_;
  assign new_n_n739_ = new_n_n181_ & new_ne2_ & new_n_n207_;
  assign new_n_n729_ = new_nk2_ & new_n_n146_ & new_n_n145_;
  assign new_n_n723_ = new_n_n147_ & new_n_n177_;
  assign new_n_n686_ = new_n_n286_ & new_nr_;
  assign new_n_n679_ = new_n_n296_ & new_n_n149_;
  assign new_nm14_ = new_n_n665_ | new_n_n667_ | new_n_n666_ | new_n_n668_;
  assign new_n_n661_ = new_ni_ & new_n_n153_ & new_nr_;
  assign new_n_n651_ = new_n_n249_ & new_n_n158_;
  assign new_n_n644_ = new_n_n260_ & new_n_n165_;
  assign new_n_n626_ = new_n_n280_ & new_nb0_;
  assign new_n_n607_ = new_n_n305_ & new_n_n161_;
  assign new_n_n600_ = new_n_n315_ & new_n_n165_;
  assign new_n_n589_ = new_ns_ & new_n_n167_ & new_nb0_;
  assign new_n_n584_ = new_n_n180_ & new_n_n168_ & new_n_n170_;
  assign new_n_n572_ = new_n_n180_ & new_n_n318_ & new_n_n172_;
  assign new_np16_ = new_n_n568_ | new_n_n566_ | new_n_n565_ | new_n_n567_ | new_n_n569_;
  assign new_n_n560_ = new_nc0_ & new_n_n182_;
  assign new_n_n555_ = new_na2_ & new_n_n207_;
  assign new_n_n553_ = new_n_n351_ & new_n_n199_ & new_n_n198_;
  assign new_np18_ = new_n_n203_ | new_nf2_;
  assign new_n_n542_ = new_ng0_ & new_n_n223_ & new_n_n210_;
  assign new_nc19_ = new_ne_ | new_nd_ | new_nc_;
  assign new_n_n536_ = new_n_n251_ & new_n_n221_ & new_n_n220_;
  assign new_n_n531_ = new_n_n225_ & new_n_n226_;
  assign new_nj20_ = new_ny1_ | new_n_n522_ | new_n_n521_;
  assign new_np20_ = new_ny1_ | new_n_n516_ | new_n_n515_;
  assign new_n_n502_ = new_n_n242_ & new_n_n244_;
  assign new_ng21_ = new_ny1_ | new_n_n500_ | new_n_n499_;
  assign new_n_n495_ = new_n_n249_ & new_ne_;
  assign new_n_n487_ = new_nd_ & new_n_n329_ & new_n_n256_;
  assign new_nt21_ = new_n_n259_ | new_n_n481_ | new_n_n480_;
  assign new_n_n473_ = new_nd_ & new_n_n329_ & new_n_n266_;
  assign new_nd22_ = new_n_n269_ | new_n_n467_ | new_n_n466_;
  assign new_n_n459_ = new_nd_ & new_n_n329_ & new_n_n276_;
  assign new_nn22_ = new_n_n279_ | new_n_n453_ | new_n_n452_;
  assign new_n_n445_ = new_nd_ & new_n_n329_ & new_n_n286_;
  assign new_nx22_ = new_n_n289_ | new_n_n439_ | new_n_n438_;
  assign new_n_n438_ = new_nd_ & new_n_n329_ & new_n_n291_;
  assign new_n_n424_ = new_nd_ & new_n_n329_ & new_n_n301_;
  assign new_nm23_ = new_n_n304_ | new_n_n418_ | new_n_n417_;
  assign new_n_n410_ = new_nd_ & new_n_n329_ & new_n_n311_;
  assign new_nw23_ = new_n_n314_ | new_n_n404_ | new_n_n403_;
  assign new_n_n396_ = new_nd_ & new_n_n329_ & new_n_n321_;
  assign new_n_n391_ = new_n_n327_ & new_ne_;
  assign new_nr24_ = new_n_n335_ | new_n_n333_ | new_n_n334_;
  assign new_nz24_ = new_nx1_ & new_n_n342_;
  assign new_n_n370_ = new_n_n363_ & new_n_n354_;
  assign new_nm25_ = new_n_n364_ | new_n_n365_;
  assign new_n_n355_ = ~new_nj25_;
  assign new_n_n346_ = ~new_nd4_;
  assign new_n_n333_ = ~new_no24_;
  assign new_n_n324_ = ~new_nx3_;
  assign new_n_n311_ = ~new_nd1_;
  assign new_n_n302_ = ~new_nu3_;
  assign new_n_n278_ = ~new_np22_;
  assign new_n_n256_ = ~new_ns0_;
  assign new_n_n247_ = ~new_nm21_;
  assign new_n_n234_ = ~new_nz2_;
  assign new_n_n225_ = ~new_ni2_;
  assign new_n_n212_ = ~new_no25_;
  assign new_n_n203_ = ~new_ne2_;
  assign new_n_n157_ = ~new_nq_;
  assign new_n_n148_ = ~new_nj_;
  assign new_n_n135_ = ~new_ny24_;
  assign new_n_n126_ = ~new_nk24_;
  assign new_n_n113_ = ~new_nm23_;
  assign new_n_n104_ = ~new_nm22_;
  assign new_n_n933_ = new_n_n124_ & new_nh2_ & new_ng2_;
  assign new_ns4_ = new_n_n13_ & new_n_n175_;
  assign new_nd5_ = new_n_n24_ & new_n_n175_;
  assign new_n_n921_ = new_n_n53_ & new_n_n52_;
  assign new_n_n915_ = new_ni2_ & new_n_n175_;
  assign new_n_n897_ = new_n_n363_ & new_no2_ & new_n_n175_;
  assign new_n_n887_ = new_n_n69_ & new_n_n70_ & new_n_n175_;
  assign new_n_n882_ = new_nx1_ & new_nr2_ & new_n_n175_;
  assign new_n_n873_ = new_n_n76_ & new_n_n235_;
  assign new_n_n863_ = new_n_n81_ & new_n_n235_;
  assign new_n_n856_ = new_n_n85_ & new_nc3_;
  assign new_n_n851_ = new_n_n87_ & new_nh_;
  assign new_n_n844_ = new_nc_ & new_n_n175_ & new_n_n91_;
  assign new_n_n826_ = new_nc_ & new_n_n175_ & new_n_n103_;
  assign new_nm7_ = new_n_n817_ | new_n_n816_ | new_n_n815_;
  assign new_n_n794_ = new_n_n126_ & new_na4_;
  assign new_n_n785_ = new_n_n335_ & new_nc4_ & new_n_n132_;
  assign new_n_n779_ = new_n_n333_ & new_nd4_ & new_n_n132_;
  assign new_n_n769_ = new_n_n337_ & new_n_n130_ & new_n_n132_;
  assign new_n_n762_ = new_n_n186_ & new_ng4_ & new_n_n132_;
  assign new_n_n754_ = new_n_n136_ & new_n_n225_;
  assign new_n_n745_ = new_n_n169_ & new_n_n139_;
  assign new_n_n737_ = new_nm2_ & new_n_n143_ & new_n_n142_;
  assign new_n_n732_ = new_nk2_ & new_n_n225_ & new_n_n145_;
  assign new_nb13_ = new_n_n722_ | new_n_n723_;
  assign new_nc14_ = new_n_n685_ | new_n_n687_ | new_n_n686_ | new_n_n688_;
  assign new_n_n680_ = new_n_n296_ & new_n_n155_;
  assign new_n_n668_ = new_n_n311_ & new_n_n155_;
  assign new_n_n659_ = new_n_n321_ & new_n_n154_;
  assign new_n_n653_ = new_ni_ & new_n_n157_ & new_nr_;
  assign new_na15_ = new_n_n641_ | new_n_n643_ | new_n_n642_ | new_n_n644_;
  assign new_n_n618_ = new_n_n290_ & new_n_n166_;
  assign new_n_n609_ = new_ns_ & new_n_n160_ & new_nb0_;
  assign new_nw15_ = new_n_n597_ | new_n_n599_ | new_n_n598_ | new_n_n600_;
  assign new_nc16_ = new_ne_ | new_n_n325_;
  assign new_n_n581_ = new_n_n180_ & new_n_n318_ & new_n_n170_;
  assign new_n_n575_ = new_n_n180_ & new_n_n171_ & new_n_n172_;
  assign new_n_n570_ = new_n_n177_ & new_n_n225_ & new_n_n180_;
  assign new_nr17_ = new_nf4_ | new_ng4_;
  assign new_n_n554_ = new_n_n201_ & new_n_n202_;
  assign new_no18_ = new_na2_ | new_n_n207_;
  assign new_nx18_ = new_ny1_ | new_n_n541_ | new_n_n540_;
  assign new_n_n537_ = new_n_n251_ & new_n_n221_ & new_n_n216_;
  assign new_nr19_ = new_nn2_ & new_nm2_ & new_nl2_;
  assign new_ny19_ = new_nx1_ | new_n_n224_ | new_n_n531_;
  assign new_n_n522_ = new_n_n231_ & new_n_n244_;
  assign new_n_n510_ = new_n_n238_ & new_n_n244_;
  assign new_ne21_ = new_ny1_ | new_n_n502_ | new_n_n501_;
  assign new_np21_ = new_n_n330_ | new_nt2_;
  assign new_nu21_ = new_n_n330_ | new_nu2_;
  assign new_n_n475_ = new_n_n263_ & new_n_n318_;
  assign new_n_n468_ = new_n_n268_ & new_n_n318_;
  assign new_nj22_ = new_n_n330_ | new_nx2_;
  assign new_no22_ = new_n_n330_ | new_ny2_;
  assign new_n_n447_ = new_n_n283_ & new_n_n318_;
  assign new_n_n440_ = new_n_n288_ & new_n_n318_;
  assign new_ni23_ = new_n_n330_ | new_nc3_;
  assign new_nn23_ = new_n_n330_ | new_nd3_;
  assign new_n_n412_ = new_n_n308_ & new_n_n318_;
  assign new_n_n405_ = new_n_n313_ & new_n_n318_;
  assign new_nc24_ = new_n_n330_ | new_ng3_;
  assign new_nj24_ = new_nn0_ | new_nl0_ | new_n_n389_;
  assign new_no24_ = new_nz3_ & new_na4_;
  assign new_n_n387_ = new_nh2_ & new_ng2_;
  assign new_nh25_ = new_no2_ | new_np2_;
  assign new_nn25_ = new_n_n361_ | new_nf0_ | new_ne0_;
  assign new_n_n358_ = ~new_nf0_;
  assign new_n_n347_ = ~new_nd25_;
  assign new_n_n332_ = ~new_nz3_;
  assign new_n_n321_ = ~new_nf1_;
  assign new_n_n314_ = ~new_nx23_;
  assign new_n_n303_ = ~new_no23_;
  assign new_n_n277_ = ~new_np3_;
  assign new_n_n266_ = ~new_nu0_;
  assign new_n_n248_ = ~new_nk21_;
  assign new_n_n233_ = ~new_ny2_;
  assign new_n_n222_ = ~new_ni25_;
  assign new_n_n215_ = ~new_nc19_;
  assign new_n_n204_ = ~new_nv16_;
  assign new_n_n178_ = ~new_nc0_;
  assign new_n_n167_ = ~new_na0_;
  assign new_n_n134_ = ~new_nw24_;
  assign new_n_n123_ = ~new_nf24_;
  assign new_n_n116_ = ~new_nq23_;
  assign new_n_n105_ = ~new_ns22_;
  assign new_n_n934_ = new_nc2_ & new_n_n124_;
  assign new_nt4_ = new_n_n14_ & new_n_n175_;
  assign new_nc5_ = new_n_n23_ & new_n_n175_;
  assign new_n_n920_ = new_n_n53_ & new_n_n54_;
  assign new_nd6_ = new_n_n914_ | new_n_n915_;
  assign new_n_n896_ = new_n_n219_ & new_no2_ & new_n_n175_;
  assign new_n_n888_ = new_n_n217_ & new_n_n70_ & new_n_n175_;
  assign new_n_n881_ = new_n_n137_ & new_nr2_ & new_n_n175_;
  assign new_n_n874_ = new_n_n76_ & new_nt2_;
  assign new_nu6_ = new_n_n861_ | new_n_n862_;
  assign new_nx6_ = new_n_n855_ | new_n_n856_;
  assign new_na7_ = new_n_n849_ | new_n_n850_;
  assign new_nd7_ = new_n_n844_ | new_n_n843_ | new_n_n842_;
  assign new_n_n825_ = new_n_n121_ & new_n_n175_ & new_n_n103_;
  assign new_n_n818_ = new_n_n108_ & new_n_n175_ & new_n_n107_;
  assign new_n_n793_ = new_nz3_ & new_ny3_ & new_n_n126_;
  assign new_n_n786_ = new_n_n332_ & new_nc4_ & new_n_n132_;
  assign new_n_n778_ = new_n_n187_ & new_nd4_ & new_n_n132_;
  assign new_n_n770_ = new_n_n336_ & new_n_n130_ & new_n_n132_;
  assign new_n_n761_ = new_n_n334_ & new_ng4_ & new_n_n132_;
  assign new_nz11_ = new_n_n754_ | new_n_n753_ | new_n_n752_;
  assign new_n_n744_ = new_n_n169_ & new_n_n141_;
  assign new_n_n738_ = new_n_n359_ & new_n_n144_ & new_n_n142_;
  assign new_n_n731_ = new_nj2_ & new_n_n225_ & new_n_n145_;
  assign new_n_n724_ = new_n_n182_ & new_nc0_;
  assign new_n_n688_ = new_n_n286_ & new_n_n155_;
  assign new_ng14_ = new_n_n677_ | new_n_n679_ | new_n_n678_ | new_n_n680_;
  assign new_n_n667_ = new_n_n311_ & new_n_n152_;
  assign new_n_n660_ = new_n_n321_ & new_n_n155_;
  assign new_nu14_ = new_n_n649_ | new_n_n651_ | new_n_n650_ | new_n_n652_;
  assign new_n_n645_ = new_ns_ & new_n_n159_ & new_n_n166_;
  assign new_n_n610_ = new_n_n300_ & new_n_n166_;
  assign new_ns15_ = new_n_n605_ | new_n_n607_ | new_n_n606_ | new_n_n608_;
  assign new_n_n601_ = new_ns_ & new_n_n162_ & new_nb0_;
  assign new_nd16_ = new_n_n224_ | new_n_n182_;
  assign new_n_n582_ = new_n_n169_ & new_n_n318_ & new_n_n170_;
  assign new_n_n574_ = new_n_n173_ & new_n_n171_ & new_n_n172_;
  assign new_no16_ = new_n_n570_ | new_n_n176_;
  assign new_nu17_ = new_nl0_ | new_n_n187_ | new_n_n188_;
  assign new_ne18_ = new_nn0_ | new_n_n341_ | new_n_n554_;
  assign new_nf18_ = new_na2_ | new_n_n203_;
  assign new_n_n541_ = new_n_n211_ & new_n_n322_;
  assign new_nh19_ = new_n_n537_ | new_ny1_;
  assign new_ns19_ = new_np2_ & new_no2_ & new_nn2_;
  assign new_n_n532_ = new_n_n223_ & new_nj2_ & new_n_n222_;
  assign new_n_n515_ = new_nf_ & new_n_n245_ & new_n_n235_;
  assign new_n_n509_ = new_nf_ & new_n_n239_ & new_nh_;
  assign new_n_n503_ = new_nf_ & new_n_n242_ & new_nh_;
  assign new_nq21_ = new_n_n485_ | new_n_n486_;
  assign new_n_n480_ = new_nd_ & new_n_n329_ & new_n_n261_;
  assign new_ny21_ = new_n_n264_ | new_n_n474_ | new_n_n473_;
  assign new_n_n469_ = new_n_n268_ & new_nx1_;
  assign new_nk22_ = new_n_n457_ | new_n_n458_;
  assign new_n_n452_ = new_nd_ & new_n_n329_ & new_n_n281_;
  assign new_ns22_ = new_n_n284_ | new_n_n446_ | new_n_n445_;
  assign new_n_n441_ = new_n_n288_ & new_nx1_;
  assign new_nj23_ = new_n_n422_ | new_n_n423_;
  assign new_n_n417_ = new_nd_ & new_n_n329_ & new_n_n306_;
  assign new_nr23_ = new_n_n309_ | new_n_n411_ | new_n_n410_;
  assign new_n_n406_ = new_n_n313_ & new_nx1_;
  assign new_nd24_ = new_n_n394_ | new_n_n395_;
  assign new_nh24_ = new_n_n330_ | new_nh3_;
  assign new_np24_ = new_n_n332_ | new_n_n335_ | new_n_n339_;
  assign new_ny24_ = new_nn0_ | new_n_n341_ | new_n_n387_;
  assign new_ni25_ = new_n_n355_ | new_n_n362_;
  assign new_n_n364_ = new_n_n360_ & new_nl2_ & new_n_n359_;
  assign new_n_n357_ = ~new_ne0_;
  assign new_n_n348_ = ~new_ne25_;
  assign new_n_n331_ = ~new_nl24_;
  assign new_n_n322_ = ~new_nk2_;
  assign new_n_n313_ = ~new_ny23_;
  assign new_n_n304_ = ~new_nn23_;
  assign new_n_n276_ = ~new_nw0_;
  assign new_n_n267_ = ~new_nn3_;
  assign new_n_n258_ = ~new_nv21_;
  assign new_n_n232_ = ~new_nx2_;
  assign new_n_n223_ = ~new_np2_;
  assign new_n_n214_ = ~new_ne19_;
  assign new_n_n205_ = ~new_ns18_;
  assign new_n_n177_ = ~new_ni3_;
  assign new_n_n168_ = ~new_nq16_;
  assign new_n_n133_ = ~new_nx24_;
  assign new_n_n124_ = ~new_nn0_;
  assign new_n_n115_ = ~new_nr23_;
  assign new_n_n106_ = ~new_nr22_;
  assign new_nn4_ = new_n_n8_ & new_n_n175_;
  assign new_nm5_ = new_n_n33_ & new_n_n175_;
  assign new_n_n930_ = new_nz1_ & new_n_n175_ & new_n_n43_;
  assign new_n_n922_ = new_n_n202_ & new_n_n51_ & new_n_n50_;
  assign new_nc6_ = new_nl0_ & new_n_n124_;
  assign new_n_n895_ = new_n_n71_ & new_no2_ & new_n_n175_;
  assign new_nl6_ = new_n_n885_ | new_n_n884_ | new_n_n883_;
  assign new_nn6_ = new_n_n875_ | new_n_n876_;
  assign new_n_n869_ = new_n_n78_ & new_n_n235_;
  assign new_n_n867_ = new_n_n79_ & new_n_n235_;
  assign new_n_n860_ = new_n_n83_ & new_na3_;
  assign new_nz6_ = new_n_n851_ | new_n_n852_;
  assign new_n_n845_ = new_n_n90_ & new_nh_;
  assign new_n_n824_ = new_n_n104_ & new_n_n175_ & new_n_n103_;
  assign new_n_n816_ = new_n_n121_ & new_n_n175_ & new_n_n109_;
  assign new_n_n808_ = new_nc_ & new_n_n175_ & new_n_n115_;
  assign new_ns7_ = new_n_n799_ | new_n_n798_ | new_n_n797_;
  assign new_ny7_ = new_n_n779_ | new_n_n777_ | new_n_n776_ | new_n_n775_ | new_n_n778_ | new_n_n780_;
  assign new_n_n771_ = new_n_n335_ & new_n_n130_ & new_n_n132_;
  assign new_nc8_ = new_n_n755_ | new_n_n756_;
  assign new_nk12_ = new_n_n750_ | new_n_n751_;
  assign new_nl12_ = new_ny1_ | new_na2_;
  assign new_no12_ = new_n_n175_ & new_na2_;
  assign new_n_n734_ = new_nj2_ & new_n_n224_ & new_n_n145_;
  assign new_n_n725_ = new_nr2_ & new_nz1_;
  assign new_n_n684_ = new_n_n291_ & new_n_n155_;
  assign new_n_n675_ = new_n_n301_ & new_n_n150_;
  assign new_nk14_ = new_n_n669_ | new_n_n671_ | new_n_n670_ | new_n_n672_;
  assign new_n_n664_ = new_n_n316_ & new_n_n155_;
  assign new_n_n655_ = new_n_n328_ & new_n_n157_;
  assign new_n_n646_ = new_n_n255_ & new_nb0_;
  assign new_nu15_ = new_n_n601_ | new_n_n603_ | new_n_n602_ | new_n_n604_;
  assign new_n_n596_ = new_n_n320_ & new_n_n165_;
  assign new_n_n593_ = new_ns_ & new_n_n164_ & new_nb0_;
  assign new_n_n587_ = new_n_n180_ & new_nq2_ & new_n_n170_;
  assign new_n_n577_ = new_n_n173_ & new_nq2_ & new_n_n172_;
  assign new_nn16_ = new_nj2_ | new_nk2_;
  assign new_n_n551_ = new_n_n204_ & new_n_n342_ & new_n_n200_;
  assign new_nr18_ = new_n_n207_ | new_ne2_ | new_nn0_;
  assign new_n_n538_ = new_n_n213_ & new_n_n360_ & new_n_n212_;
  assign new_no19_ = new_no2_ & new_nn2_ & new_nm2_;
  assign new_n_n533_ = new_n_n222_ & new_n_n360_;
  assign new_nh21_ = new_n_n251_ & new_n_n329_;
  assign new_n_n493_ = new_ni3_ & new_nx1_;
  assign new_n_n477_ = new_n_n263_ & new_n_n262_;
  assign new_n_n470_ = new_n_n268_ & new_n_n267_;
  assign new_n_n437_ = new_nq3_ & new_nx1_;
  assign new_n_n430_ = new_nr3_ & new_nx1_;
  assign new_n_n407_ = new_n_n313_ & new_n_n312_;
  assign new_n_n395_ = new_nw3_ & new_nx1_;
  assign new_n_n385_ = new_n_n346_ & new_n_n349_ & new_n_n347_;
  assign new_n_n376_ = new_n_n354_ & new_nf4_ & new_n_n350_;
  assign new_n_n330_ = ~new_nl21_;
  assign new_n_n319_ = ~new_nc24_;
  assign new_n_n297_ = ~new_nt3_;
  assign new_n_n286_ = ~new_ny0_;
  assign new_n_n231_ = ~new_nw2_;
  assign new_n_n220_ = ~new_nc16_;
  assign new_n_n209_ = ~new_nw18_;
  assign new_n_n198_ = ~new_nk18_;
  assign new_n_n187_ = ~new_nj17_;
  assign new_n_n132_ = ~new_nh17_;
  assign new_n_n121_ = ~new_nh21_;
  assign new_n_n110_ = ~new_nb23_;
  assign new_n_n99_ = ~new_nd22_;
  assign new_n_n8_ = ~new_nq13_;
  assign new_nm4_ = new_n_n7_ & new_n_n175_;
  assign new_nn5_ = new_n_n34_ & new_n_n175_;
  assign new_n_n931_ = new_n_n325_ & new_n_n42_ & new_n_n41_;
  assign new_ny5_ = new_n_n920_ | new_n_n921_;
  assign new_nb6_ = new_n_n124_ & new_nh2_;
  assign new_n_n894_ = new_n_n363_ & new_n_n68_ & new_n_n175_;
  assign new_n_n886_ = new_n_n71_ & new_n_n70_ & new_n_n175_;
  assign new_n_n876_ = new_n_n75_ & new_ns2_;
  assign new_n_n870_ = new_n_n78_ & new_nv2_;
  assign new_ns6_ = new_n_n865_ | new_n_n866_;
  assign new_nv6_ = new_n_n859_ | new_n_n860_;
  assign new_n_n852_ = new_n_n87_ & new_ne3_;
  assign new_n_n846_ = new_n_n90_ & new_nh3_;
  assign new_nk7_ = new_n_n823_ | new_n_n822_ | new_n_n821_;
  assign new_n_n817_ = new_nc_ & new_n_n175_ & new_n_n109_;
  assign new_n_n807_ = new_n_n121_ & new_n_n175_ & new_n_n115_;
  assign new_n_n800_ = new_n_n120_ & new_n_n175_ & new_n_n119_;
  assign new_n_n780_ = new_n_n335_ & new_nd4_ & new_n_n132_;
  assign new_n_n772_ = new_n_n337_ & new_ne4_ & new_n_n132_;
  assign new_n_n756_ = new_n_n135_ & new_nh4_;
  assign new_nj12_ = new_nk2_ | new_nj2_ | new_na2_;
  assign new_nn12_ = new_n_n748_ | new_n_n746_ | new_n_n745_ | new_n_n747_ | new_n_n749_ | new_n_n744_ | new_n_n743_ | new_n_n742_ | new_n_n741_;
  assign new_n_n741_ = new_n_n140_ & new_n_n141_;
  assign new_n_n733_ = new_n_n173_ & new_n_n224_ & new_n_n145_;
  assign new_n_n726_ = new_nz1_ & new_nc0_;
  assign new_n_n683_ = new_n_n291_ & new_n_n148_;
  assign new_n_n676_ = new_n_n301_ & new_n_n155_;
  assign new_n_n672_ = new_n_n306_ & new_n_n155_;
  assign new_no14_ = new_n_n661_ | new_n_n663_ | new_n_n662_ | new_n_n664_;
  assign new_n_n654_ = new_n_n328_ & new_n_n156_;
  assign new_n_n647_ = new_n_n255_ & new_n_n159_;
  assign new_n_n604_ = new_n_n310_ & new_n_n165_;
  assign new_ny15_ = new_n_n593_ | new_n_n595_ | new_n_n594_ | new_n_n596_;
  assign new_na16_ = new_n_n589_ | new_n_n591_ | new_n_n590_ | new_n_n592_;
  assign new_n_n588_ = new_n_n169_ & new_nq2_ & new_n_n170_;
  assign new_n_n576_ = new_nq12_ & new_n_n171_ & new_n_n172_;
  assign new_nm16_ = new_n_n182_ & new_n_n177_;
  assign new_n_n550_ = new_n_n206_ & new_n_n342_ & new_n_n200_;
  assign new_n_n547_ = new_n_n205_ & new_n_n206_;
  assign new_n_n545_ = new_n_n209_ & new_n_n323_;
  assign new_nq19_ = new_n_n536_ | new_n_n218_;
  assign new_nx19_ = new_n_n532_ | new_n_n533_;
  assign new_ni21_ = new_n_n498_ | new_n_n497_ | new_n_n496_;
  assign new_nm21_ = new_n_n492_ | new_n_n493_;
  assign new_n_n476_ = new_n_n263_ & new_nx1_;
  assign new_nc22_ = new_n_n470_ | new_n_n469_ | new_n_n468_;
  assign new_n_n436_ = new_n_n323_ & new_n_n322_ & new_nq3_;
  assign new_ne23_ = new_n_n429_ | new_n_n430_;
  assign new_n_n413_ = new_n_n308_ & new_nx1_;
  assign new_n_n389_ = new_nz3_ & new_ny3_;
  assign new_n_n384_ = new_n_n351_ & new_n_n349_ & new_n_n347_;
  assign new_n_n377_ = new_n_n353_ & new_n_n354_ & new_n_n350_;
  assign new_n_n329_ = ~new_ne_;
  assign new_n_n320_ = ~new_nv1_;
  assign new_n_n296_ = ~new_na1_;
  assign new_n_n287_ = ~new_nr3_;
  assign new_n_n230_ = ~new_nv2_;
  assign new_n_n221_ = ~new_nc_;
  assign new_n_n199_ = ~new_nj18_;
  assign new_n_n197_ = ~new_nf4_;
  assign new_n_n188_ = ~new_nk17_;
  assign new_n_n131_ = ~new_nv24_;
  assign new_n_n122_ = ~new_ng24_;
  assign new_n_n109_ = ~new_nc23_;
  assign new_n_n100_ = ~new_nc22_;
  assign new_nw4_ = new_n_n17_ & new_n_n175_;
  assign new_nh5_ = new_n_n28_ & new_n_n175_;
  assign new_no5_ = new_n_n35_ & new_n_n175_;
  assign new_nw5_ = new_n_n928_ | new_n_n926_ | new_n_n925_ | new_n_n924_ | new_n_n927_ | new_n_n929_;
  assign new_nx5_ = new_n_n922_ | new_n_n923_;
  assign new_n_n916_ = new_n_n124_ & new_n_n61_ & new_n_n60_;
  assign new_n_n893_ = new_n_n219_ & new_n_n68_ & new_n_n175_;
  assign new_n_n884_ = new_n_n72_ & new_nx1_;
  assign new_n_n878_ = new_n_n137_ & new_n_n73_ & new_n_n175_;
  assign new_nq6_ = new_n_n869_ | new_n_n870_;
  assign new_n_n866_ = new_n_n80_ & new_nx2_;
  assign new_nw6_ = new_n_n857_ | new_n_n858_;
  assign new_n_n854_ = new_n_n86_ & new_nd3_;
  assign new_nc7_ = new_n_n845_ | new_n_n846_;
  assign new_n_n823_ = new_nc_ & new_n_n175_ & new_n_n105_;
  assign new_nn7_ = new_n_n814_ | new_n_n813_ | new_n_n812_;
  assign new_n_n809_ = new_n_n114_ & new_n_n175_ & new_n_n113_;
  assign new_n_n801_ = new_n_n121_ & new_n_n175_ & new_n_n119_;
  assign new_nu7_ = new_n_n795_ | new_n_n796_;
  assign new_n_n788_ = new_n_n335_ & new_n_n127_ & new_n_n132_;
  assign new_n_n758_ = new_n_n334_ & new_n_n133_ & new_n_n132_;
  assign new_ni12_ = new_n_n169_ | new_ny1_;
  assign new_n_n749_ = new_n_n325_ & new_n_n138_;
  assign new_n_n740_ = new_nd0_ & new_n_n203_ & new_nf2_;
  assign new_nw12_ = new_n_n734_ | new_n_n732_ | new_n_n731_ | new_n_n733_ | new_n_n735_ | new_n_n730_ | new_n_n729_ | new_n_n728_ | new_n_n727_;
  assign new_na13_ = new_n_n726_ | new_n_n725_ | new_n_n724_;
  assign new_n_n685_ = new_ni_ & new_n_n157_ & new_n_n156_;
  assign new_ni14_ = new_n_n673_ | new_n_n675_ | new_n_n674_ | new_n_n676_;
  assign new_n_n671_ = new_n_n306_ & new_n_n151_;
  assign new_n_n662_ = new_n_n316_ & new_n_n156_;
  assign new_ns14_ = new_n_n653_ | new_n_n655_ | new_n_n654_ | new_n_n656_;
  assign new_n_n648_ = new_n_n255_ & new_n_n165_;
  assign new_n_n606_ = new_n_n305_ & new_n_n166_;
  assign new_n_n597_ = new_ns_ & new_n_n163_ & new_nb0_;
  assign new_n_n592_ = new_n_n327_ & new_n_n165_;
  assign new_n_n585_ = new_n_n169_ & new_n_n168_ & new_n_n170_;
  assign new_n_n579_ = new_nq12_ & new_nq2_ & new_n_n172_;
  assign new_nl16_ = new_n_n323_ & new_n_n322_;
  assign new_nh18_ = new_n_n552_ | new_n_n551_ | new_n_n550_;
  assign new_n_n548_ = new_n_n205_ & new_n_n204_;
  assign new_n_n544_ = new_n_n325_ & new_nj2_ & new_nw18_;
  assign new_nb19_ = new_n_n363_ & new_nx1_ & new_n_n215_;
  assign new_n_n534_ = new_n_n225_ & new_n_n224_ & new_n_n226_;
  assign new_n_n500_ = new_n_n243_ & new_n_n244_;
  assign new_nl21_ = new_n_n329_ & new_n_n251_ & new_nc_;
  assign new_n_n489_ = new_n_n253_ & new_n_n318_;
  assign new_n_n482_ = new_n_n258_ & new_n_n318_;
  assign new_ny22_ = new_n_n330_ | new_na3_;
  assign new_nd23_ = new_n_n330_ | new_nb3_;
  assign new_n_n419_ = new_n_n303_ & new_n_n318_;
  assign new_ns24_ = new_n_n346_ & new_nc4_ & new_nb4_;
  assign new_n_n386_ = new_n_n351_ & new_n_n346_;
  assign new_n_n378_ = new_nk0_ & new_nf4_ & new_ng4_;
  assign new_n_n310_ = ~new_nt1_;
  assign new_n_n299_ = ~new_ni23_;
  assign new_n_n288_ = ~new_nz22_;
  assign new_n_n229_ = ~new_nu2_;
  assign new_n_n211_ = ~new_nz18_;
  assign new_n_n200_ = ~new_ni18_;
  assign new_n_n130_ = ~new_nr24_;
  assign new_n_n119_ = ~new_nb24_;
  assign new_n_n112_ = ~new_ng23_;
  assign new_n_n101_ = ~new_ni22_;
  assign new_nx4_ = new_n_n18_ & new_n_n175_;
  assign new_ng5_ = new_n_n27_ & new_n_n175_;
  assign new_np5_ = new_n_n36_ & new_n_n175_;
  assign new_nv5_ = new_n_n44_ & new_n_n175_;
  assign new_n_n923_ = new_n_n49_ & new_n_n48_ & new_n_n127_;
  assign new_n_n917_ = new_n_n124_ & new_n_n59_ & new_n_n58_;
  assign new_n_n892_ = new_n_n71_ & new_n_n68_ & new_n_n175_;
  assign new_n_n885_ = new_n_n72_ & new_n_n224_;
  assign new_n_n877_ = new_n_n74_ & new_n_n73_ & new_n_n175_;
  assign new_n_n871_ = new_n_n77_ & new_n_n235_;
  assign new_n_n865_ = new_n_n80_ & new_n_n235_;
  assign new_n_n859_ = new_n_n83_ & new_nh_;
  assign new_n_n853_ = new_n_n86_ & new_nh_;
  assign new_n_n847_ = new_n_n89_ & new_nh_;
  assign new_n_n822_ = new_n_n121_ & new_n_n175_ & new_n_n105_;
  assign new_n_n815_ = new_n_n110_ & new_n_n175_ & new_n_n109_;
  assign new_np7_ = new_n_n808_ | new_n_n807_ | new_n_n806_;
  assign new_n_n802_ = new_nc_ & new_n_n175_ & new_n_n119_;
  assign new_n_n796_ = new_n_n125_ & new_nz3_;
  assign new_n_n789_ = new_n_n332_ & new_n_n127_ & new_n_n132_;
  assign new_n_n757_ = new_n_n134_ & new_n_n133_ & new_n_n132_;
  assign new_nc12_ = new_nq2_ & new_nr2_;
  assign new_n_n748_ = new_n_n325_ & new_n_n139_;
  assign new_np12_ = new_n_n739_ | new_n_n740_;
  assign new_n_n735_ = new_nk2_ & new_n_n224_ & new_n_n145_;
  assign new_nz12_ = new_n_n562_ | new_n_n225_;
  assign new_ne14_ = new_n_n681_ | new_n_n683_ | new_n_n682_ | new_n_n684_;
  assign new_n_n677_ = new_ni_ & new_n_n149_ & new_nr_;
  assign new_n_n670_ = new_n_n306_ & new_n_n156_;
  assign new_n_n663_ = new_n_n316_ & new_n_n153_;
  assign new_n_n656_ = new_n_n328_ & new_n_n155_;
  assign new_ny14_ = new_n_n645_ | new_n_n647_ | new_n_n646_ | new_n_n648_;
  assign new_n_n605_ = new_ns_ & new_n_n161_ & new_nb0_;
  assign new_n_n598_ = new_n_n315_ & new_n_n166_;
  assign new_n_n591_ = new_n_n327_ & new_n_n167_;
  assign new_n_n586_ = new_n_n173_ & new_nq2_ & new_n_n170_;
  assign new_n_n578_ = new_n_n180_ & new_nq2_ & new_n_n172_;
  assign new_nj16_ = new_ni2_ & new_n_n175_ & new_n_n325_;
  assign new_n_n552_ = new_nh0_ & new_n_n342_ & new_n_n200_;
  assign new_n_n549_ = new_n_n205_ & new_nh0_;
  assign new_nw18_ = new_n_n542_ | new_n_n543_;
  assign new_na19_ = new_nd_ | new_nc_ | new_n_n214_;
  assign new_nn19_ = new_nl2_ & new_nm2_;
  assign new_n_n499_ = new_nf_ & new_n_n245_ & new_nh_;
  assign new_nk21_ = new_n_n330_ | new_ns2_;
  assign new_no21_ = new_n_n254_ | new_n_n488_ | new_n_n487_;
  assign new_n_n483_ = new_n_n258_ & new_nx1_;
  assign new_nz22_ = new_n_n436_ | new_n_n437_;
  assign new_n_n431_ = new_nd_ & new_n_n329_ & new_n_n296_;
  assign new_nh23_ = new_n_n299_ | new_n_n425_ | new_n_n424_;
  assign new_nb25_ = new_n_n344_ | new_n_n345_ | new_n_n386_;
  assign new_nc25_ = new_n_n382_ | new_n_n384_ | new_n_n383_ | new_n_n385_;
  assign new_n_n379_ = new_n_n353_ & new_nk0_ & new_ng4_;
  assign new_n_n309_ = ~new_ns23_;
  assign new_n_n300_ = ~new_nr1_;
  assign new_n_n298_ = ~new_nj23_;
  assign new_n_n219_ = ~new_no19_;
  assign new_n_n210_ = ~new_nl25_;
  assign new_n_n201_ = ~new_nd2_;
  assign new_n_n129_ = ~new_np24_;
  assign new_n_n120_ = ~new_na24_;
  assign new_n_n111_ = ~new_nh23_;
  assign new_n_n102_ = ~new_nh22_;
  assign new_ni5_ = new_n_n29_ & new_n_n175_;
  assign new_nt5_ = new_n_n932_ | new_nn0_;
  assign new_n_n925_ = new_n_n336_ & new_n_n46_ & new_n_n132_;
  assign new_na6_ = new_n_n57_ | new_n_n917_ | new_n_n916_;
  assign new_ng6_ = new_n_n908_ | new_n_n909_;
  assign new_n_n901_ = new_n_n71_ & new_nn2_ & new_n_n175_;
  assign new_n_n848_ = new_n_n89_ & new_ng3_;
  assign new_n_n838_ = new_nc_ & new_n_n175_ & new_n_n95_;
  assign new_ni7_ = new_n_n829_ | new_n_n828_ | new_n_n827_;
  assign new_n_n720_ = new_ni3_ & new_n_n225_;
  assign new_n_n711_ = new_n_n256_ & new_n_n149_;
  assign new_n_n702_ = new_n_n266_ & new_nr_;
  assign new_n_n693_ = new_ni_ & new_n_n153_ & new_n_n156_;
  assign new_nc15_ = new_n_n637_ | new_n_n639_ | new_n_n638_ | new_n_n640_;
  assign new_n_n632_ = new_n_n275_ & new_n_n165_;
  assign new_n_n623_ = new_n_n285_ & new_n_n167_;
  assign new_n_n614_ = new_n_n295_ & new_n_n166_;
  assign new_n_n566_ = new_n_n178_ & new_n_n325_ & new_nd0_;
  assign new_n_n559_ = new_n_n183_ & new_nh0_;
  assign new_ne17_ = new_n_n349_ & new_nd4_ & new_nc4_;
  assign new_ny17_ = new_n_n192_ & new_n_n191_ & new_n_n190_;
  assign new_nk18_ = new_n_n201_ | new_n_n202_ | new_nk0_;
  assign new_n_n521_ = new_nf_ & new_n_n235_ & new_n_n232_;
  assign new_n_n514_ = new_n_n236_ & new_n_n244_;
  assign new_na21_ = new_ny1_ | new_n_n506_ | new_n_n505_;
  assign new_n_n496_ = new_n_n247_ & new_n_n318_;
  assign new_n_n490_ = new_n_n253_ & new_nx1_;
  assign new_np22_ = new_n_n450_ | new_n_n451_;
  assign new_nu22_ = new_n_n443_ | new_n_n444_;
  assign new_n_n434_ = new_n_n293_ & new_nx1_;
  assign new_n_n427_ = new_n_n298_ & new_nx1_;
  assign new_n_n420_ = new_n_n303_ & new_nx1_;
  assign new_nt24_ = new_ny3_ & new_nz3_;
  assign new_nd25_ = new_n_n348_ | new_n_n381_ | new_n_n380_;
  assign new_n_n373_ = new_n_n363_ & new_n_n352_;
  assign new_nl25_ = new_n_n362_ | new_n_n356_ | new_n_n366_;
  assign new_n_n359_ = ~new_nm2_;
  assign new_n_n293_ = ~new_ne23_;
  assign new_n_n282_ = ~new_nq3_;
  assign new_n_n271_ = ~new_nv0_;
  assign new_n_n260_ = ~new_nj1_;
  assign new_n_n249_ = ~new_nh1_;
  assign new_n_n194_ = ~new_nd18_;
  assign new_n_n183_ = ~new_nx16_;
  assign new_n_n172_ = ~new_no16_;
  assign new_n_n161_ = ~new_nw_;
  assign new_n_n150_ = ~new_nl_;
  assign new_n_n139_ = ~new_no12_;
  assign new_n_n4_ = ~new_nj12_;
  assign new_nj5_ = new_n_n30_ & new_n_n175_;
  assign new_ns5_ = new_n_n536_ | new_ny1_;
  assign new_n_n924_ = new_n_n47_ & new_n_n46_ & new_n_n132_;
  assign new_n_n918_ = new_n_n124_ & new_n_n203_ & new_n_n56_;
  assign new_n_n909_ = new_n_n363_ & new_n_n175_ & new_n_n64_;
  assign new_n_n902_ = new_n_n66_ & new_nn2_ & new_n_n175_;
  assign new_ny6_ = new_n_n853_ | new_n_n854_;
  assign new_n_n837_ = new_n_n121_ & new_n_n175_ & new_n_n95_;
  assign new_n_n830_ = new_n_n100_ & new_n_n175_ & new_n_n99_;
  assign new_n_n719_ = new_ni3_ & new_nq2_;
  assign new_n_n712_ = new_n_n256_ & new_n_n155_;
  assign new_n_n701_ = new_ni_ & new_n_n151_ & new_n_n156_;
  assign new_n_n694_ = new_n_n276_ & new_nr_;
  assign new_n_n640_ = new_n_n265_ & new_n_n165_;
  assign new_ng15_ = new_n_n629_ | new_n_n631_ | new_n_n630_ | new_n_n632_;
  assign new_n_n622_ = new_n_n285_ & new_nb0_;
  assign new_n_n615_ = new_n_n295_ & new_n_n159_;
  assign new_n_n565_ = new_n_n325_ & new_n_n224_ & new_nd0_;
  assign new_nt16_ = new_n_n559_ | new_n_n558_ | new_n_n557_;
  assign new_ng17_ = new_n_n186_ | new_n_n187_ | new_n_n188_;
  assign new_nx17_ = new_nn0_ | new_n_n189_;
  assign new_nu18_ = new_ny1_ | new_n_n545_ | new_n_n544_;
  assign new_n_n528_ = new_n_n228_ & new_n_n244_;
  assign new_n_n513_ = new_nf_ & new_n_n237_ & new_nh_;
  assign new_n_n507_ = new_nf_ & new_n_n240_ & new_nh_;
  assign new_nj21_ = new_n_n248_ | new_n_n495_ | new_n_n494_;
  assign new_n_n491_ = new_n_n253_ & new_n_n252_;
  assign new_n_n451_ = new_no3_ & new_nx1_;
  assign new_nt22_ = new_n_n330_ | new_nz2_;
  assign new_n_n433_ = new_n_n293_ & new_n_n318_;
  assign new_n_n428_ = new_n_n298_ & new_n_n297_;
  assign new_n_n414_ = new_n_n308_ & new_n_n307_;
  assign new_nk24_ = new_nn0_ | new_nl0_ | new_n_n388_;
  assign new_n_n381_ = new_ni0_ & new_n_n349_;
  assign new_n_n374_ = new_nl2_ & new_n_n351_;
  assign new_n_n366_ = new_n_n360_ & new_n_n358_ & new_n_n357_;
  assign new_n_n360_ = ~new_no2_;
  assign new_n_n292_ = ~new_ns3_;
  assign new_n_n283_ = ~new_nu22_;
  assign new_n_n270_ = ~new_nl1_;
  assign new_n_n261_ = ~new_nt0_;
  assign new_n_n239_ = ~new_nd3_;
  assign new_n_n193_ = ~new_nb2_;
  assign new_n_n184_ = ~new_na25_;
  assign new_n_n171_ = ~new_nm16_;
  assign new_n_n162_ = ~new_nx_;
  assign new_n_n149_ = ~new_nk_;
  assign new_n_n140_ = ~new_nr12_;
  assign new_n_n5_ = ~new_ni12_;
  assign new_nk5_ = new_n_n31_ & new_n_n175_;
  assign new_nu5_ = new_n_n40_ | new_n_n931_ | new_n_n930_;
  assign new_n_n927_ = new_n_n47_ & new_nb2_ & new_n_n132_;
  assign new_n_n919_ = new_n_n124_ & new_n_n55_ & new_n_n59_;
  assign new_n_n911_ = new_n_n63_ & new_nk2_;
  assign new_n_n903_ = new_n_n363_ & new_nn2_ & new_n_n175_;
  assign new_n_n861_ = new_n_n82_ & new_n_n235_;
  assign new_n_n839_ = new_n_n94_ & new_n_n175_ & new_n_n93_;
  assign new_n_n831_ = new_n_n121_ & new_n_n175_ & new_n_n99_;
  assign new_n_n718_ = new_nd0_ & new_ni2_ & new_nr2_;
  assign new_n_n709_ = new_ni_ & new_n_n149_ & new_n_n156_;
  assign new_n_n704_ = new_n_n266_ & new_n_n155_;
  assign new_n_n695_ = new_n_n276_ & new_n_n153_;
  assign new_n_n682_ = new_n_n291_ & new_n_n156_;
  assign new_n_n639_ = new_n_n265_ & new_n_n161_;
  assign new_n_n630_ = new_n_n275_ & new_nb0_;
  assign new_nk15_ = new_n_n621_ | new_n_n623_ | new_n_n622_ | new_n_n624_;
  assign new_n_n616_ = new_n_n295_ & new_n_n165_;
  assign new_n_n603_ = new_n_n310_ & new_n_n162_;
  assign new_n_n594_ = new_n_n320_ & new_n_n166_;
  assign new_nq16_ = new_n_n182_ & new_ni3_;
  assign new_n_n557_ = new_n_n183_ & new_n_n206_;
  assign new_nc17_ = new_ny3_ & new_nb2_ & new_n_n185_;
  assign new_nw17_ = new_n_n196_ | new_n_n332_ | new_n_n335_;
  assign new_ni18_ = new_n_n208_ & new_nh4_;
  assign new_n_n546_ = new_nh4_ & new_n_n208_;
  assign new_n_n527_ = new_nf_ & new_n_n235_ & new_n_n229_;
  assign new_n_n520_ = new_n_n232_ & new_n_n244_;
  assign new_n_n508_ = new_n_n239_ & new_n_n244_;
  assign new_n_n498_ = new_n_n247_ & new_n_n246_;
  assign new_nn21_ = new_n_n491_ | new_n_n490_ | new_n_n489_;
  assign new_n_n464_ = new_n_n323_ & new_n_n322_ & new_nm3_;
  assign new_n_n457_ = new_n_n323_ & new_n_n322_ & new_nn3_;
  assign new_nb23_ = new_n_n435_ | new_n_n434_ | new_n_n433_;
  assign new_ng23_ = new_n_n428_ | new_n_n427_ | new_n_n426_;
  assign new_nv23_ = new_n_n407_ | new_n_n406_ | new_n_n405_;
  assign new_n_n394_ = new_n_n323_ & new_n_n322_ & new_nw3_;
  assign new_n_n383_ = new_n_n346_ & new_ni0_ & new_n_n347_;
  assign new_n_n375_ = new_n_n352_ & new_n_n351_;
  assign new_n_n350_ = ~new_ng4_;
  assign new_n_n339_ = ~new_nm24_;
  assign new_n_n295_ = ~new_nq1_;
  assign new_n_n284_ = ~new_nt22_;
  assign new_n_n269_ = ~new_ne22_;
  assign new_n_n251_ = ~new_nd_;
  assign new_n_n240_ = ~new_ne3_;
  assign new_n_n196_ = ~new_na4_;
  assign new_n_n185_ = ~new_nr17_;
  assign new_n_n170_ = ~new_nr16_;
  assign new_n_n159_ = ~new_nu_;
  assign new_n_n152_ = ~new_nn_;
  assign new_n_n141_ = ~new_np12_;
  assign new_n_n6_ = ~new_nl12_;
  assign new_nl5_ = new_n_n32_ & new_n_n175_;
  assign new_n_n932_ = new_ni2_ & new_n_n325_ & new_n_n39_;
  assign new_n_n926_ = new_n_n45_ & new_n_n46_ & new_n_n132_;
  assign new_nz5_ = new_n_n918_ | new_n_n919_;
  assign new_n_n910_ = new_n_n63_ & new_n_n325_;
  assign new_ni6_ = new_n_n902_ | new_n_n900_ | new_n_n899_ | new_n_n898_ | new_n_n901_ | new_n_n903_;
  assign new_n_n868_ = new_n_n79_ & new_nw2_;
  assign new_nf7_ = new_n_n838_ | new_n_n837_ | new_n_n836_;
  assign new_n_n832_ = new_nc_ & new_n_n175_ & new_n_n99_;
  assign new_n_n717_ = new_nd0_ & new_nr2_ & new_ni3_;
  assign new_n_n710_ = new_n_n256_ & new_nr_;
  assign new_n_n703_ = new_n_n266_ & new_n_n151_;
  assign new_n_n696_ = new_n_n276_ & new_n_n155_;
  assign new_n_n674_ = new_n_n301_ & new_n_n156_;
  assign new_n_n638_ = new_n_n265_ & new_nb0_;
  assign new_n_n631_ = new_n_n275_ & new_n_n163_;
  assign new_n_n624_ = new_n_n285_ & new_n_n165_;
  assign new_no15_ = new_n_n613_ | new_n_n615_ | new_n_n614_ | new_n_n616_;
  assign new_n_n602_ = new_n_n310_ & new_n_n166_;
  assign new_n_n595_ = new_n_n320_ & new_n_n164_;
  assign new_nr16_ = new_n_n564_ | new_n_n179_;
  assign new_n_n558_ = new_n_n183_ & new_n_n204_;
  assign new_nd17_ = new_nb4_ & new_na4_ & new_nz3_;
  assign new_nv17_ = new_nc2_ | new_n_n193_ | new_nn0_;
  assign new_nj18_ = new_ni0_ | new_nj0_;
  assign new_ns18_ = new_n_n546_ | new_na2_;
  assign new_nf20_ = new_ny1_ | new_n_n526_ | new_n_n525_;
  assign new_nl20_ = new_ny1_ | new_n_n520_ | new_n_n519_;
  assign new_ns20_ = new_ny1_ | new_n_n514_ | new_n_n513_;
  assign new_n_n497_ = new_n_n247_ & new_nx1_;
  assign new_n_n492_ = new_n_n323_ & new_n_n322_ & new_ni3_;
  assign new_nh22_ = new_n_n463_ | new_n_n462_ | new_n_n461_;
  assign new_n_n458_ = new_nn3_ & new_nx1_;
  assign new_n_n435_ = new_n_n293_ & new_n_n292_;
  assign new_n_n429_ = new_n_n323_ & new_n_n322_ & new_nr3_;
  assign new_n_n401_ = new_n_n323_ & new_n_n322_ & new_nv3_;
  assign new_na24_ = new_n_n400_ | new_n_n399_ | new_n_n398_;
  assign new_n_n382_ = new_n_n351_ & new_ni0_ & new_n_n347_;
  assign new_nf25_ = new_n_n373_ | new_n_n375_ | new_n_n374_ | new_n_n362_;
  assign new_n_n349_ = ~new_ne4_;
  assign new_n_n340_ = ~new_nu24_;
  assign new_n_n294_ = ~new_nd23_;
  assign new_n_n285_ = ~new_no1_;
  assign new_n_n259_ = ~new_nu21_;
  assign new_n_n250_ = ~new_nr0_;
  assign new_n_n241_ = ~new_nf3_;
  assign new_n_n195_ = ~new_nb4_;
  assign new_n_n186_ = ~new_ni17_;
  assign new_n_n169_ = ~new_nq12_;
  assign new_n_n160_ = ~new_nv_;
  assign new_n_n151_ = ~new_nm_;
  assign new_n_n142_ = ~new_nh25_;
  assign new_n_n7_ = ~new_nm13_;
  assign new_n_n937_ = new_n_n221_ & new_n_n1_ & new_n_n0_;
  assign new_nq4_ = new_n_n11_ & new_n_n175_;
  assign new_nb5_ = new_n_n22_ & new_n_n175_;
  assign new_n_n912_ = new_n_n62_ & new_n_n325_;
  assign new_n_n904_ = new_nm2_ & new_n_n71_ & new_n_n65_;
  assign new_no6_ = new_n_n873_ | new_n_n874_;
  assign new_n_n841_ = new_nc_ & new_n_n175_ & new_n_n93_;
  assign new_nh7_ = new_n_n832_ | new_n_n831_ | new_n_n830_;
  assign new_nm13_ = new_n_n713_ | new_n_n715_ | new_n_n714_ | new_n_n716_;
  assign new_n_n708_ = new_n_n261_ & new_n_n155_;
  assign new_n_n699_ = new_n_n271_ & new_n_n152_;
  assign new_n_n690_ = new_n_n281_ & new_nr_;
  assign new_n_n666_ = new_n_n311_ & new_n_n156_;
  assign new_n_n637_ = new_ns_ & new_n_n161_ & new_n_n166_;
  assign new_ni15_ = new_n_n625_ | new_n_n627_ | new_n_n626_ | new_n_n628_;
  assign new_n_n620_ = new_n_n290_ & new_n_n165_;
  assign new_n_n611_ = new_n_n300_ & new_n_n160_;
  assign new_nf16_ = new_ny1_ | new_nz1_;
  assign new_nh16_ = new_n_n578_ | new_n_n576_ | new_n_n575_ | new_n_n577_ | new_n_n579_ | new_n_n574_ | new_n_n573_ | new_n_n572_ | new_n_n571_;
  assign new_n_n564_ = new_ni3_ & new_n_n225_ & new_n_n180_;
  assign new_nw16_ = new_nd2_ & new_nl0_ & new_n_n354_;
  assign new_nj17_ = new_nd4_ & new_nc4_ & new_nb4_;
  assign new_nd18_ = new_n_n197_ & new_n_n350_;
  assign new_n_n540_ = new_n_n325_ & new_nk2_ & new_nz18_;
  assign new_nj19_ = new_nm2_ & new_nn2_;
  assign new_n_n535_ = new_nx1_ & new_n_n224_;
  assign new_n_n526_ = new_n_n229_ & new_n_n244_;
  assign new_nn20_ = new_ny1_ | new_n_n518_ | new_n_n517_;
  assign new_n_n511_ = new_nf_ & new_n_n238_ & new_nh_;
  assign new_n_n504_ = new_n_n241_ & new_n_n244_;
  assign new_n_n486_ = new_nj3_ & new_nx1_;
  assign new_n_n479_ = new_nk3_ & new_nx1_;
  assign new_n_n472_ = new_nl3_ & new_nx1_;
  assign new_n_n465_ = new_nm3_ & new_nx1_;
  assign new_n_n463_ = new_n_n273_ & new_n_n272_;
  assign new_n_n456_ = new_n_n278_ & new_n_n277_;
  assign new_n_n449_ = new_n_n283_ & new_n_n282_;
  assign new_n_n442_ = new_n_n288_ & new_n_n287_;
  assign new_n_n423_ = new_ns3_ & new_nx1_;
  assign new_n_n416_ = new_nt3_ & new_nx1_;
  assign new_n_n409_ = new_nu3_ & new_nx1_;
  assign new_n_n402_ = new_nv3_ & new_nx1_;
  assign new_n_n400_ = new_n_n317_ & new_n_n324_;
  assign new_n_n393_ = new_nk2_ & new_n_n325_;
  assign new_nm24_ = new_nc4_ & new_nb4_ & new_na4_;
  assign new_nx24_ = new_n_n338_ | new_n_n339_ | new_n_n340_;
  assign new_nj25_ = new_n_n369_ | new_n_n368_ | new_n_n367_;
  assign new_n_n363_ = ~new_nl2_;
  assign new_n_n352_ = ~new_ni0_;
  assign new_n_n341_ = ~new_nb_;
  assign new_n_n338_ = ~new_nt24_;
  assign new_n_n327_ = ~new_nw1_;
  assign new_n_n316_ = ~new_ne1_;
  assign new_n_n305_ = ~new_ns1_;
  assign new_n_n289_ = ~new_ny22_;
  assign new_n_n275_ = ~new_nm1_;
  assign new_n_n264_ = ~new_nz21_;
  assign new_n_n253_ = ~new_nq21_;
  assign new_n_n242_ = ~new_ng3_;
  assign new_n_n228_ = ~new_nt2_;
  assign new_n_n217_ = ~new_nn19_;
  assign new_n_n206_ = ~new_nw16_;
  assign new_n_n190_ = ~new_nb18_;
  assign new_n_n179_ = ~new_ns16_;
  assign new_n_n176_ = ~new_np16_;
  assign new_n_n165_ = ~new_ns_;
  assign new_n_n154_ = ~new_np_;
  assign new_n_n143_ = ~new_ng25_;
  assign new_n_n118_ = ~new_nv23_;
  assign new_n_n107_ = ~new_nx22_;
  assign new_n_n0_ = ~new_nz11_;
  assign new_nj4_ = new_n_n937_ | new_ny1_;
  assign new_nr4_ = new_n_n12_ & new_n_n175_;
  assign new_na5_ = new_n_n21_ & new_n_n175_;
  assign new_nf6_ = new_n_n910_ | new_n_n911_;
  assign new_n_n905_ = new_nl2_ & new_n_n71_ & new_n_n65_;
  assign new_nm6_ = new_n_n881_ | new_n_n879_ | new_n_n878_ | new_n_n877_ | new_n_n880_ | new_n_n882_;
  assign new_n_n840_ = new_n_n121_ & new_n_n175_ & new_n_n93_;
  assign new_n_n833_ = new_n_n98_ & new_n_n175_ & new_n_n97_;
  assign new_n_n716_ = new_n_n250_ & new_n_n155_;
  assign new_ns13_ = new_n_n705_ | new_n_n707_ | new_n_n706_ | new_n_n708_;
  assign new_n_n698_ = new_n_n271_ & new_nr_;
  assign new_n_n691_ = new_n_n281_ & new_n_n154_;
  assign new_n_n658_ = new_n_n321_ & new_n_n156_;
  assign new_ne15_ = new_n_n633_ | new_n_n635_ | new_n_n634_ | new_n_n636_;
  assign new_n_n629_ = new_ns_ & new_n_n163_ & new_n_n166_;
  assign new_n_n619_ = new_n_n290_ & new_n_n158_;
  assign new_n_n612_ = new_n_n300_ & new_n_n165_;
  assign new_ng16_ = new_n_n587_ | new_n_n585_ | new_n_n584_ | new_n_n586_ | new_n_n588_ | new_n_n583_ | new_n_n582_ | new_n_n581_ | new_n_n580_;
  assign new_n_n580_ = new_n_n173_ & new_n_n318_ & new_n_n170_;
  assign new_ns16_ = new_n_n563_ | new_n_n561_ | new_n_n560_ | new_n_n562_ | new_n_n225_;
  assign new_nv16_ = new_n_n352_ & new_n_n353_;
  assign new_nk17_ = new_n_n350_ & new_n_n197_ & new_n_n349_;
  assign new_nb18_ = new_ne4_ | new_n_n346_ | new_n_n344_;
  assign new_nz18_ = new_n_n538_ | new_n_n539_;
  assign new_ni19_ = new_nm2_ | new_n_n325_ | new_ne_;
  assign new_nd20_ = new_ny1_ | new_n_n528_ | new_n_n527_;
  assign new_n_n525_ = new_nf_ & new_n_n235_ & new_n_n230_;
  assign new_n_n519_ = new_nf_ & new_n_n235_ & new_n_n233_;
  assign new_nw20_ = new_ny1_ | new_n_n510_ | new_n_n509_;
  assign new_nc21_ = new_ny1_ | new_n_n504_ | new_n_n503_;
  assign new_n_n485_ = new_n_n323_ & new_n_n322_ & new_nj3_;
  assign new_nv21_ = new_n_n478_ | new_n_n479_;
  assign new_n_n471_ = new_n_n323_ & new_n_n322_ & new_nl3_;
  assign new_nf22_ = new_n_n464_ | new_n_n465_;
  assign new_n_n462_ = new_n_n273_ & new_nx1_;
  assign new_nm22_ = new_n_n456_ | new_n_n455_ | new_n_n454_;
  assign new_n_n448_ = new_n_n283_ & new_nx1_;
  assign new_nw22_ = new_n_n442_ | new_n_n441_ | new_n_n440_;
  assign new_n_n422_ = new_n_n323_ & new_n_n322_ & new_ns3_;
  assign new_no23_ = new_n_n415_ | new_n_n416_;
  assign new_n_n408_ = new_n_n323_ & new_n_n322_ & new_nu3_;
  assign new_ny23_ = new_n_n401_ | new_n_n402_;
  assign new_n_n399_ = new_n_n317_ & new_nx1_;
  assign new_nf24_ = new_n_n324_ | new_n_n393_ | new_n_n392_;
  assign new_nn24_ = new_n_n332_ | new_n_n335_ | new_n_n331_;
  assign new_nw24_ = new_ng4_ & new_nf4_ & new_ne4_;
  assign new_n_n369_ = new_n_n361_ & new_nl2_ & new_n_n359_;
  assign new_no25_ = new_n_n362_ | new_nm2_ | new_n_n363_;
  assign new_n_n351_ = ~new_nh0_;
  assign new_n_n342_ = ~new_na2_;
  assign new_n_n337_ = ~new_nq24_;
  assign new_n_n328_ = ~new_ng1_;
  assign new_n_n315_ = ~new_nu1_;
  assign new_n_n306_ = ~new_nc1_;
  assign new_n_n279_ = ~new_no22_;
  assign new_n_n274_ = ~new_nj22_;
  assign new_n_n265_ = ~new_nk1_;
  assign new_n_n252_ = ~new_nk3_;
  assign new_n_n243_ = ~new_nh3_;
  assign new_n_n238_ = ~new_nc3_;
  assign new_n_n216_ = ~new_ni19_;
  assign new_n_n207_ = ~new_nf2_;
  assign new_n_n189_ = ~new_nc2_;
  assign new_n_n180_ = ~new_nl16_;
  assign new_n_n175_ = ~new_ny1_;
  assign new_n_n166_ = ~new_nb0_;
  assign new_n_n153_ = ~new_no_;
  assign new_n_n144_ = ~new_nf25_;
  assign new_n_n117_ = ~new_nw23_;
  assign new_n_n108_ = ~new_nw22_;
  assign new_n_n1_ = ~new_ny11_;
  assign new_n_n936_ = new_n_n5_ & new_n_n4_ & new_n_n3_;
  assign new_no4_ = new_n_n9_ & new_n_n175_;
  assign new_nz4_ = new_n_n20_ & new_n_n175_;
  assign new_ne6_ = new_n_n912_ | new_n_n913_;
  assign new_n_n906_ = new_nl2_ & new_n_n359_ & new_n_n65_;
  assign new_n_n891_ = new_n_n217_ & new_np2_ & new_n_n175_;
  assign new_n_n715_ = new_n_n250_ & new_n_n148_;
  assign new_n_n706_ = new_n_n261_ & new_nr_;
  assign new_nw13_ = new_n_n697_ | new_n_n699_ | new_n_n698_ | new_n_n700_;
  assign new_n_n692_ = new_n_n281_ & new_n_n155_;
  assign new_n_n650_ = new_n_n249_ & new_nb0_;
  assign new_n_n636_ = new_n_n270_ & new_n_n165_;
  assign new_n_n627_ = new_n_n280_ & new_n_n164_;
  assign new_n_n621_ = new_ns_ & new_n_n167_ & new_n_n166_;
  assign new_nq15_ = new_n_n609_ | new_n_n611_ | new_n_n610_ | new_n_n612_;
  assign new_n_n571_ = new_n_n173_ & new_n_n318_ & new_n_n172_;
  assign new_n_n567_ = new_n_n325_ & new_n_n224_ & new_n_n182_;
  assign new_n_n563_ = new_n_n224_ & new_n_n181_;
  assign new_n_n556_ = new_na2_ & new_n_n203_;
  assign new_nh17_ = new_nl0_ | new_nn0_;
  assign new_na18_ = new_n_n195_ | new_n_n196_ | new_n_n332_;
  assign new_n_n539_ = new_np2_ & new_n_n360_ & new_n_n212_;
  assign new_nv19_ = new_nx19_ | new_ni2_;
  assign new_n_n529_ = new_nf_ & new_n_n235_ & new_n_n228_;
  assign new_nh20_ = new_ny1_ | new_n_n524_ | new_n_n523_;
  assign new_n_n517_ = new_nf_ & new_n_n235_ & new_n_n234_;
  assign new_nu20_ = new_ny1_ | new_n_n512_ | new_n_n511_;
  assign new_n_n505_ = new_nf_ & new_n_n241_ & new_nh_;
  assign new_ns21_ = new_n_n484_ | new_n_n483_ | new_n_n482_;
  assign new_nx21_ = new_n_n477_ | new_n_n476_ | new_n_n475_;
  assign new_nz21_ = new_n_n330_ | new_nv2_;
  assign new_ne22_ = new_n_n330_ | new_nw2_;
  assign new_n_n461_ = new_n_n273_ & new_n_n318_;
  assign new_n_n454_ = new_n_n278_ & new_n_n318_;
  assign new_n_n450_ = new_n_n323_ & new_n_n322_ & new_no3_;
  assign new_n_n443_ = new_n_n323_ & new_n_n322_ & new_np3_;
  assign new_nc23_ = new_n_n294_ | new_n_n432_ | new_n_n431_;
  assign new_nl23_ = new_n_n421_ | new_n_n420_ | new_n_n419_;
  assign new_nq23_ = new_n_n414_ | new_n_n413_ | new_n_n412_;
  assign new_ns23_ = new_n_n330_ | new_ne3_;
  assign new_nx23_ = new_n_n330_ | new_nf3_;
  assign new_n_n398_ = new_n_n317_ & new_n_n318_;
  assign new_ng24_ = new_n_n326_ | new_n_n391_ | new_n_n390_;
  assign new_n_n388_ = new_ny3_ & new_nz3_ & new_na4_;
  assign new_nv24_ = new_n_n335_ | new_n_n336_ | new_n_n337_;
  assign new_n_n380_ = new_n_n353_ & new_nf4_;
  assign new_n_n372_ = new_n_n354_ & new_n_n353_;
  assign new_n_n368_ = new_no2_ & new_nl2_ & new_n_n359_;
  assign new_n_n361_ = ~new_ng0_;
  assign new_n_n354_ = ~new_nk0_;
  assign new_n_n343_ = ~new_nb25_;
  assign new_n_n336_ = ~new_nd17_;
  assign new_n_n325_ = ~new_nx1_;
  assign new_n_n318_ = ~new_nn16_;
  assign new_n_n307_ = ~new_nv3_;
  assign new_n_n291_ = ~new_nz0_;
  assign new_n_n280_ = ~new_nn1_;
  assign new_n_n273_ = ~new_nk22_;
  assign new_n_n262_ = ~new_nm3_;
  assign new_n_n255_ = ~new_ni1_;
  assign new_n_n244_ = ~new_nf_;
  assign new_n_n237_ = ~new_nb3_;
  assign new_n_n226_ = ~new_nx19_;
  assign new_n_n208_ = ~new_ny16_;
  assign new_n_n192_ = ~new_nz17_;
  assign new_n_n181_ = ~new_nd0_;
  assign new_n_n174_ = ~new_nj16_;
  assign new_n_n163_ = ~new_ny_;
  assign new_n_n156_ = ~new_nr_;
  assign new_n_n145_ = ~new_nb13_;
  assign new_n_n138_ = ~new_nm0_;
  assign new_n_n127_ = ~new_nw17_;
  assign new_n_n2_ = ~new_nn12_;
  assign new_nk4_ = new_n_n2_ | new_n_n936_ | new_n_n935_;
  assign new_np4_ = new_n_n10_ & new_n_n175_;
  assign new_ny4_ = new_n_n19_ & new_n_n175_;
  assign new_n_n913_ = new_n_n62_ & new_nj2_;
  assign new_n_n907_ = new_n_n363_ & new_nm2_ & new_n_n65_;
  assign new_n_n899_ = new_n_n66_ & new_n_n67_ & new_n_n175_;
  assign new_n_n714_ = new_n_n250_ & new_nr_;
  assign new_n_n707_ = new_n_n261_ & new_n_n150_;
  assign new_n_n700_ = new_n_n271_ & new_n_n155_;
  assign new_na14_ = new_n_n689_ | new_n_n691_ | new_n_n690_ | new_n_n692_;
  assign new_n_n642_ = new_n_n260_ & new_nb0_;
  assign new_n_n635_ = new_n_n270_ & new_n_n162_;
  assign new_n_n628_ = new_n_n280_ & new_n_n165_;
  assign new_nm15_ = new_n_n617_ | new_n_n619_ | new_n_n618_ | new_n_n620_;
  assign new_n_n613_ = new_ns_ & new_n_n159_ & new_nb0_;
  assign new_ni16_ = new_n_n182_ | new_n_n224_ | new_n_n174_;
  assign new_n_n568_ = new_n_n178_ & new_n_n325_ & new_n_n182_;
  assign new_n_n562_ = new_n_n182_ & new_n_n224_;
  assign new_nx16_ = new_n_n556_ | new_n_n555_ | new_n_n546_;
  assign new_ni17_ = new_na4_ & new_nz3_ & new_ny3_;
  assign new_nz17_ = new_n_n335_ | new_n_n193_ | new_n_n194_;
  assign new_nl19_ = new_n_n536_ | new_n_n217_;
  assign new_nw19_ = new_ny1_ | new_n_n535_ | new_n_n534_;
  assign new_n_n530_ = new_n_n227_ & new_n_n244_;
  assign new_n_n524_ = new_n_n230_ & new_n_n244_;
  assign new_n_n518_ = new_n_n233_ & new_n_n244_;
  assign new_n_n512_ = new_n_n237_ & new_n_n244_;
  assign new_n_n506_ = new_n_n240_ & new_n_n244_;
  assign new_n_n484_ = new_n_n258_ & new_n_n257_;
  assign new_n_n478_ = new_n_n323_ & new_n_n322_ & new_nk3_;
  assign new_na22_ = new_n_n471_ | new_n_n472_;
  assign new_n_n466_ = new_nd_ & new_n_n329_ & new_n_n271_;
  assign new_ni22_ = new_n_n274_ | new_n_n460_ | new_n_n459_;
  assign new_n_n455_ = new_n_n278_ & new_nx1_;
  assign new_nr22_ = new_n_n449_ | new_n_n448_ | new_n_n447_;
  assign new_n_n444_ = new_np3_ & new_nx1_;
  assign new_n_n426_ = new_n_n298_ & new_n_n318_;
  assign new_n_n421_ = new_n_n303_ & new_n_n302_;
  assign new_n_n415_ = new_n_n323_ & new_n_n322_ & new_nt3_;
  assign new_nt23_ = new_n_n408_ | new_n_n409_;
  assign new_n_n403_ = new_nd_ & new_n_n329_ & new_n_n316_;
  assign new_nb24_ = new_n_n319_ | new_n_n397_ | new_n_n396_;
  assign new_n_n392_ = new_nj2_ & new_n_n325_;
  assign new_nl24_ = new_na4_ & new_nb4_;
  assign new_nu24_ = new_nf4_ & new_ne4_ & new_n_n346_;
  assign new_ne25_ = new_n_n376_ | new_n_n378_ | new_n_n377_ | new_n_n379_;
  assign new_ng25_ = new_n_n370_ | new_n_n372_ | new_n_n371_ | new_nn2_;
  assign new_n_n367_ = new_np2_ & new_nl2_ & new_n_n359_;
  assign new_n_n362_ = ~new_nn2_;
  assign new_n_n353_ = ~new_nj0_;
  assign new_n_n344_ = ~new_nc4_;
  assign new_n_n335_ = ~new_ny3_;
  assign new_n_n326_ = ~new_nh24_;
  assign new_n_n317_ = ~new_nd24_;
  assign new_n_n308_ = ~new_nt23_;
  assign new_n_n290_ = ~new_np1_;
  assign new_n_n281_ = ~new_nx0_;
  assign new_n_n272_ = ~new_no3_;
  assign new_n_n263_ = ~new_na22_;
  assign new_n_n254_ = ~new_np21_;
  assign new_n_n245_ = ~new_ng_;
  assign new_n_n236_ = ~new_na3_;
  assign new_n_n227_ = ~new_ns2_;
  assign new_n_n218_ = ~new_nr19_;
  assign new_n_n191_ = ~new_na18_;
  assign new_n_n182_ = ~new_nr2_;
  assign new_n_n173_ = ~new_nz12_;
  assign new_n_n164_ = ~new_nz_;
  assign new_n_n155_ = ~new_ni_;
  assign new_n_n146_ = ~new_na13_;
  assign new_n_n137_ = ~new_nc12_;
  assign new_n_n128_ = ~new_nn24_;
  assign new_n_n3_ = ~new_nk12_;
  assign new_n_n93_ = ~new_no21_;
  assign new_n_n82_ = ~new_np20_;
  assign new_n_n71_ = ~new_na19_;
  assign new_n_n60_ = ~new_nq18_;
  assign new_n_n49_ = ~new_nu17_;
  assign new_n_n94_ = ~new_nn21_;
  assign new_n_n81_ = ~new_nn20_;
  assign new_n_n72_ = ~new_nw19_;
  assign new_n_n59_ = ~new_ng18_;
  assign new_n_n50_ = ~new_ny17_;
  assign new_n_n95_ = ~new_nt21_;
  assign new_n_n80_ = ~new_nl20_;
  assign new_n_n69_ = ~new_ns19_;
  assign new_n_n62_ = ~new_nu18_;
  assign new_n_n51_ = ~new_nx17_;
  assign new_n_n96_ = ~new_ns21_;
  assign new_n_n79_ = ~new_nj20_;
  assign new_n_n70_ = ~new_nu19_;
  assign new_n_n61_ = ~new_np18_;
  assign new_n_n52_ = ~new_nh2_;
  assign new_ni4_ = ~new_nz24_;
  assign new_n_n835_ = new_nc_ & new_n_n175_ & new_n_n97_;
  assign new_nj7_ = new_n_n826_ | new_n_n825_ | new_n_n824_;
  assign new_n_n705_ = new_ni_ & new_n_n150_ & new_n_n156_;
  assign new_ny13_ = new_n_n693_ | new_n_n695_ | new_n_n694_ | new_n_n696_;
  assign new_n_n617_ = new_ns_ & new_n_n158_ & new_nb0_;
  assign new_n_n97_ = ~new_ny21_;
  assign new_n_n42_ = ~new_nf16_;
  assign new_n_n31_ = ~new_nm15_;
  assign new_n_n20_ = ~new_no14_;
  assign new_n_n9_ = ~new_ns13_;
  assign new_n_n834_ = new_n_n121_ & new_n_n175_ & new_n_n97_;
  assign new_n_n827_ = new_n_n102_ & new_n_n175_ & new_n_n101_;
  assign new_nu13_ = new_n_n701_ | new_n_n703_ | new_n_n702_ | new_n_n704_;
  assign new_n_n697_ = new_ni_ & new_n_n152_ & new_n_n156_;
  assign new_n_n625_ = new_ns_ & new_n_n164_ & new_n_n166_;
  assign new_n_n98_ = ~new_nx21_;
  assign new_n_n41_ = ~new_ng16_;
  assign new_n_n32_ = ~new_no15_;
  assign new_n_n19_ = ~new_nm14_;
  assign new_n_n10_ = ~new_nu13_;
  assign new_n_n908_ = new_n_n71_ & new_n_n175_ & new_n_n64_;
  assign new_n_n836_ = new_n_n96_ & new_n_n175_ & new_n_n95_;
  assign new_n_n828_ = new_n_n121_ & new_n_n175_ & new_n_n101_;
  assign new_nc13_ = new_n_n720_ | new_n_n718_ | new_n_n717_ | new_n_n719_ | new_n_n721_;
  assign new_nq13_ = new_n_n709_ | new_n_n711_ | new_n_n710_ | new_n_n712_;
  assign new_n_n633_ = new_ns_ & new_n_n162_ & new_n_n166_;
  assign new_n_n40_ = ~new_ni16_;
  assign new_n_n29_ = ~new_ni15_;
  assign new_n_n22_ = ~new_ns14_;
  assign new_n_n11_ = ~new_nw13_;
  assign new_n_n900_ = new_n_n363_ & new_n_n67_ & new_n_n175_;
  assign new_ng7_ = new_n_n835_ | new_n_n834_ | new_n_n833_;
  assign new_n_n829_ = new_nc_ & new_n_n175_ & new_n_n101_;
  assign new_n_n721_ = new_nq2_ & new_ni2_;
  assign new_n_n713_ = new_ni_ & new_n_n148_ & new_n_n156_;
  assign new_n_n641_ = new_ns_ & new_n_n160_ & new_n_n166_;
  assign new_n_n39_ = ~new_nd16_;
  assign new_n_n30_ = ~new_nk15_;
  assign new_n_n21_ = ~new_nq14_;
  assign new_n_n12_ = ~new_ny13_;
  assign new_nk6_ = new_n_n890_ | new_n_n888_ | new_n_n887_ | new_n_n886_ | new_n_n889_ | new_n_n891_;
  assign new_n_n821_ = new_n_n106_ & new_n_n175_ & new_n_n105_;
  assign new_n_n813_ = new_n_n121_ & new_n_n175_ & new_n_n111_;
  assign new_n_n805_ = new_nc_ & new_n_n175_ & new_n_n117_;
  assign new_nt7_ = new_n_n335_ & new_n_n124_ & new_n_n202_;
  assign new_n_n736_ = new_n_n144_ & new_n_n143_ & new_n_n142_;
  assign new_n_n727_ = new_n_n173_ & new_n_n146_ & new_n_n145_;
  assign new_n_n649_ = new_ns_ & new_n_n158_ & new_n_n166_;
  assign new_n_n68_ = ~new_nq19_;
  assign new_n_n57_ = ~new_nr18_;
  assign new_n_n46_ = ~new_ng17_;
  assign new_n_n35_ = ~new_nu15_;
  assign new_n_n24_ = ~new_ny14_;
  assign new_n_n13_ = ~new_na14_;
  assign new_n_n883_ = new_n_n72_ & new_n_n74_;
  assign new_nl7_ = new_n_n820_ | new_n_n819_ | new_n_n818_;
  assign new_n_n814_ = new_nc_ & new_n_n175_ & new_n_n111_;
  assign new_n_n804_ = new_n_n121_ & new_n_n175_ & new_n_n117_;
  assign new_n_n797_ = new_n_n123_ & new_n_n175_ & new_n_n122_;
  assign new_nr12_ = new_n_n175_ & new_n_n342_;
  assign new_n_n728_ = new_nj2_ & new_n_n146_ & new_n_n145_;
  assign new_n_n657_ = new_ni_ & new_n_n154_ & new_nr_;
  assign new_n_n67_ = ~new_nl19_;
  assign new_n_n58_ = ~new_no18_;
  assign new_n_n45_ = ~new_nc17_;
  assign new_n_n36_ = ~new_nw15_;
  assign new_n_n23_ = ~new_nu14_;
  assign new_n_n14_ = ~new_nc14_;
  assign new_n_n875_ = new_n_n75_ & new_n_n235_;
  assign new_n_n820_ = new_nc_ & new_n_n175_ & new_n_n107_;
  assign new_no7_ = new_n_n811_ | new_n_n810_ | new_n_n809_;
  assign new_n_n806_ = new_n_n116_ & new_n_n175_ & new_n_n115_;
  assign new_n_n798_ = new_n_n121_ & new_n_n175_ & new_n_n122_;
  assign new_n_n751_ = new_ni2_ & new_nr2_;
  assign new_n_n742_ = new_n_n140_ & new_n_n139_;
  assign new_n_n665_ = new_ni_ & new_n_n152_ & new_nr_;
  assign new_n_n88_ = ~new_nc21_;
  assign new_n_n77_ = ~new_nf20_;
  assign new_n_n44_ = ~new_nt16_;
  assign new_n_n33_ = ~new_nq15_;
  assign new_n_n26_ = ~new_nc15_;
  assign new_n_n15_ = ~new_ne14_;
  assign new_nr6_ = new_n_n867_ | new_n_n868_;
  assign new_n_n819_ = new_n_n121_ & new_n_n175_ & new_n_n107_;
  assign new_n_n812_ = new_n_n112_ & new_n_n175_ & new_n_n111_;
  assign new_nq7_ = new_n_n805_ | new_n_n804_ | new_n_n803_;
  assign new_n_n799_ = new_nc_ & new_n_n175_ & new_n_n122_;
  assign new_n_n750_ = new_ni2_ & new_nq2_;
  assign new_n_n743_ = new_n_n140_ & new_n_n138_;
  assign new_n_n673_ = new_ni_ & new_n_n150_ & new_nr_;
  assign new_n_n87_ = ~new_na21_;
  assign new_n_n78_ = ~new_nh20_;
  assign new_n_n43_ = ~new_nh16_;
  assign new_n_n34_ = ~new_ns15_;
  assign new_n_n25_ = ~new_na15_;
  assign new_n_n16_ = ~new_ng14_;
  assign new_n_n862_ = new_n_n82_ & new_nz2_;
  assign new_nw7_ = new_n_n791_ | new_n_n789_ | new_n_n788_ | new_n_n787_ | new_n_n790_ | new_n_n792_;
  assign new_n_n783_ = new_n_n332_ & new_n_n128_ & new_n_n132_;
  assign new_n_n774_ = new_n_n335_ & new_ne4_ & new_n_n132_;
  assign new_n_n764_ = new_n_n339_ & new_n_n131_ & new_n_n132_;
  assign new_n_n763_ = new_n_n340_ & new_n_n131_ & new_n_n132_;
  assign new_ny11_ = new_nd_ | new_ne_;
  assign new_n_n681_ = new_ni_ & new_n_n148_ & new_nr_;
  assign new_n_n89_ = ~new_ne21_;
  assign new_n_n86_ = ~new_ny20_;
  assign new_n_n75_ = ~new_na20_;
  assign new_n_n64_ = ~new_nb19_;
  assign new_n_n53_ = ~new_ne18_;
  assign new_n_n28_ = ~new_ng15_;
  assign new_n_n17_ = ~new_ni14_;
  assign new_n_n855_ = new_n_n85_ & new_nh_;
  assign new_n_n792_ = new_n_n332_ & new_nb4_ & new_n_n132_;
  assign new_n_n784_ = new_n_n339_ & new_nc4_ & new_n_n132_;
  assign new_n_n773_ = new_n_n336_ & new_ne4_ & new_n_n132_;
  assign new_n_n765_ = new_n_n338_ & new_n_n131_ & new_n_n132_;
  assign new_nb8_ = new_n_n761_ | new_n_n759_ | new_n_n758_ | new_n_n757_ | new_n_n760_ | new_n_n762_;
  assign new_n_n755_ = new_nd2_ & new_nl0_ & new_n_n135_;
  assign new_n_n689_ = new_ni_ & new_n_n154_ & new_n_n156_;
  assign new_n_n90_ = ~new_ng21_;
  assign new_n_n85_ = ~new_nw20_;
  assign new_n_n76_ = ~new_nd20_;
  assign new_n_n63_ = ~new_nx18_;
  assign new_n_n54_ = ~new_ng2_;
  assign new_n_n27_ = ~new_ne15_;
  assign new_n_n18_ = ~new_nk14_;
  assign new_nb7_ = new_n_n847_ | new_n_n848_;
  assign new_n_n791_ = new_n_n335_ & new_nb4_ & new_n_n132_;
  assign new_n_n781_ = new_n_n339_ & new_n_n128_ & new_n_n132_;
  assign new_n_n775_ = new_n_n187_ & new_n_n129_ & new_n_n132_;
  assign new_n_n766_ = new_n_n340_ & new_nf4_ & new_n_n132_;
  assign new_n_n91_ = ~new_nj21_;
  assign new_n_n84_ = ~new_nu20_;
  assign new_n_n73_ = ~new_ny19_;
  assign new_n_n66_ = ~new_nj19_;
  assign new_n_n55_ = ~new_nf18_;
  assign new_n_n48_ = ~new_nv17_;
  assign new_n_n37_ = ~new_ny15_;
  assign new_ne7_ = new_n_n841_ | new_n_n840_ | new_n_n839_;
  assign new_n_n790_ = new_n_n331_ & new_nb4_ & new_n_n132_;
  assign new_n_n782_ = new_n_n335_ & new_n_n128_ & new_n_n132_;
  assign new_nz7_ = new_n_n773_ | new_n_n771_ | new_n_n770_ | new_n_n769_ | new_n_n772_ | new_n_n774_;
  assign new_n_n767_ = new_n_n339_ & new_nf4_ & new_n_n132_;
  assign new_n_n92_ = ~new_ni21_;
  assign new_n_n83_ = ~new_ns20_;
  assign new_n_n74_ = ~new_nv19_;
  assign new_n_n65_ = ~new_nh19_;
  assign new_n_n56_ = ~new_nh18_;
  assign new_n_n47_ = ~new_ne17_;
  assign new_n_n38_ = ~new_na16_;
endmodule


