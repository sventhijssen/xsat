// Benchmark "spla" written by ABC on Sat Apr 29 10:30:21 2023

module spla ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
    f0, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15,
    f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26, f27, f28, f29,
    f30, f31, f32, f33, f34, f35, f36, f37, f38, f39, f40, f41, f42, f43,
    f44, f45  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15;
  output f0, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15,
    f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26, f27, f28, f29,
    f30, f31, f32, f33, f34, f35, f36, f37, f38, f39, f40, f41, f42, f43,
    f44, f45;
  assign f0 = x0 & (~x1 | (~x7 & ~x4 & ~x6 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & ~x14 & ~x3 & ~x2 & x5));
  assign f1 = x2 ? ~x0 : (x0 & (~x1 | (~x4 & ~x6 & ~x8 & ~x9 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & ~x14 & ~x3 & x5 & x7)));
  assign f2 = x0 & x5 & x1 & ~x2 & ~x3 & ~x14 & ~x15 & ~x13 & ~x12 & ~x11 & ~x10 & ~x9 & ~x8 & ~x4 & ~x6;
  assign f3 = ~x3 & ~x4 & ((~x5 & ~x2 & ~x0 & x1 & (x7 | (~x11 & ~x12 & ((~x13 & (x8 ? (~x15 & ~x14 & (~x9 | ~x10)) : ((x9 | x10) & (x15 ^ x14)))) | (~x8 & x13 & ~x15 & ~x14 & (x9 | x10)))))) | (x0 & ~x1));
  assign f4 = ~x3 & x4 & ((~x5 & ~x2 & ~x0 & x1 & (x7 | (~x11 & ~x12 & ((~x8 & (x9 | x10) & (x13 ? (~x15 & ~x14) : (x15 ^ x14))) | (~x13 & ~x15 & ~x14 & x8 & (x9 ^ x10)))))) | (x0 & ~x1));
  assign f5 = ~x3 & ((~x2 & ((x4 & ((((x12 & ~x13) | (~x15 & x14)) & ((~x0 & ~x5 & ((x7 & ~x10 & x6 & ~x11 & (x9 ^ x8)) | (~x1 & (~x7 | ~x6)))) | (~x1 & x5 & (x7 | (x10 & x6 & ~x11))))) | (x6 & ((~x0 & ~x5 & ((~x12 & ~x11 & ((~x13 & ((~x15 & ((x9 & ~x10 & (x8 ? (~x14 & x1) : x14)) | (x10 & ((~x7 & ~x8 & x14) | (~x9 & x8 & ~x14 & x1))))) | (~x8 & x15 & ~x14 & x1 & (x9 | x10)))) | (~x8 & x13 & ~x15 & ~x14 & x1 & (x9 | x10)))) | (x7 & x1))) | (x12 & x14 & ~x10 & x11 & ~x1 & x5 & (x13 ^ x15)))))) | (~x0 & ~x1 & ~x4 & ((x5 & ((x12 & ~x13) | (~x15 & x14)) & ((~x9 & (x8 ? (~x10 & ~x11) : (~x6 & (x10 ^ x11)))) | ~x7 | (~x10 & ~x11 & (x6 | (x9 & ~x8))))) | (x10 & ~x11 & ~x5 & (x7 ^ x6)))))) | (x0 & ~x1 & x5 & x4));
  assign f6 = ~x4 & ~x3 & ((~x2 & x6 & ~x5 & ~x0 & x1 & (x7 | (~x11 & ~x12 & ((~x13 & (x8 ? (~x15 & ~x14 & (~x9 | ~x10)) : ((x9 | x10) & (x15 ^ x14)))) | (~x8 & x13 & ~x15 & ~x14 & (x9 | x10)))))) | (x5 & x0 & ~x1));
  assign f7 = ~x1 & ~x3 & ~x2 & ~x0 & ((((x13 & x12) | (x15 & x14)) & (((~x4 ^ ~x5) & (~x7 | (~x10 & ~x11 & (x8 ^ x9)))) | (x5 & (x4 ? (x7 | (x6 & ~x10 & x11)) : ((~x8 & ~x9 & ~x6 & (~x10 ^ ~x11)) | (x6 & ~x10 & ~x11)))) | (~x6 & x4 & ~x5))) | (x6 & ((x12 & x14 & x10 & ~x11 & x4 & x5 & (x13 ^ x15)) | (~x7 & ~x10 & x11 & ~x4 & ~x5))) | (x11 & ~x4 & ~x5 & x7 & ~x6 & ~x10));
  assign f8 = x3 & ~x1 & ~x0;
  assign f9 = (~x7 | ((x8 | ((x9 | ((~x6 | x5) & (x6 | x10 | x11 | x4))) & (x4 | ((~x10 | ~x11) & (~x6 | (~x10 & ~x11)))))) & ((~x10 & ~x11) | ((~x6 | x5 | ~x4) & (~x8 | ~x5 | x4))) & (~x9 | ((~x8 | (x6 ? x5 : (x10 | x4))) & (x4 | (~x11 & (~x10 | ~x5))))))) & (~x5 | (((~x14 ^ ~x15) | (x12 ^ x13)) & (x7 | ~x4 | ((x12 | (x14 & (x15 | ~x11))) & (~x11 | (~x10 & (x13 | (x14 & x15)))) & x6 & (x11 | (x10 & (~x15 | ~x13))))))) & (~x4 | (~x14 ^ ~x15) | (x12 ^ x13)) & (x5 | x4 | (((x6 & x7) | (x10 & ~x11)) & (~x9 | x10) & (x6 | x7))) & ~x0 & ~x2 & ~x3 & ~x1;
  assign f10 = ~x3 & ((~x2 & ((~x0 & ((((x15 & ~x14) | (~x12 & x13)) & ((x7 & x4 & (x5 ? ~x1 : ~x6)) | (~x1 & x5 & ~x4 & ((~x9 & (x8 ? (~x10 & ~x11) : (~x6 & (~x10 ^ ~x11)))) | ~x7 | (~x10 & ~x11 & (x6 | (x9 & ~x8))))))) | (~x5 & ((x7 & ((~x6 & x1 & x4) | (~x9 & x8 & x6 & ~x1 & ~x4))) | (~x6 & ~x12 & ~x11 & x4 & ((~x13 & ((~x15 & x1 & ((x9 & (x8 ? (~x14 & ~x10) : x14)) | (x10 & ((~x8 & x14) | (~x9 & x8 & ~x14))))) | (~x8 & x15 & ~x14 & (x9 | x10)))) | (~x8 & x13 & ~x15 & ~x14 & (x9 | x10)))))) | (x6 & ~x1 & x5 & x4 & ((x15 & ((x12 & ~x14 & (x13 ? (~x10 & x11) : (x10 & ~x11))) | (~x12 & x13 & x14 & ~x10 & x11))) | (x14 & x10 & ~x11 & ~x12 & x13 & ~x15))))) | (~x1 & ~x5 & x4 & (~x7 | (~x10 & ~x11 & (x9 ^ x8))) & ((x15 & ~x14) | (~x12 & x13))))) | (x0 & ~x1 & ~x5 & x4));
  assign f11 = ~x5 & ~x4 & ~x3 & ((x0 & ~x1) | (~x6 & ~x2 & ~x0 & x1 & (x7 | (~x11 & ~x12 & ((~x13 & (x8 ? (~x15 & ~x14 & (~x9 | ~x10)) : ((x9 | x10) & (x15 ^ x14)))) | (~x8 & x13 & ~x15 & ~x14 & (x9 | x10)))))));
  assign f12 = ~x1 & ~x3 & ~x2 & ~x0 & (x5 ? ((((~x13 & ~x12) | (~x15 & ~x14)) & (x4 ? x7 : ((~x8 & (x9 ? (~x10 & ~x11) : (~x6 & (~x10 ^ ~x11)))) | ~x7 | (~x10 & ~x11 & (x6 | (x8 & ~x9)))))) | (x6 & x4 & ((~x15 & ((~x13 & x10 & ~x11 & (x12 ^ x14)) | (x13 & x12 & ~x14 & ~x10 & x11))) | (x14 & ~x10 & x11 & ~x13 & ~x12 & x15)))) : ((x4 & ((~x13 & ~x12) | (~x15 & ~x14)) & ((~x10 & ~x11 & (x8 ^ x9)) | ~x7 | ~x6)) | (x7 & ~x8 & x9 & x6 & ~x4)));
  assign f13 = ~x1 & ~x3 & ~x2 & ~x0 & x6 & (x7 ? (x4 & x5) : (~x4 & ~x5 & (~x10 ^ ~x11)));
  assign f14 = x4 & ~x0 & ~x2 & ~x3 & ~x6 & ~x5 & ~x1 & ~x7;
  assign f15 = ~x1 & ~x10 & ~x11 & ~x3 & ~x2 & ~x0 & x7 & x6 & (x5 ? ~x4 : (x4 & (~x8 ^ ~x9)));
  assign f16 = ~x1 & ~x4 & ~x6 & ~x3 & ~x2 & ~x0 & x5 & x7 & ((~x8 & (x9 ? (~x10 & ~x11) : (~x10 ^ ~x11))) | (~x10 & ~x11 & x8 & ~x9));
  assign f17 = x4 & x7 & ~x0 & ~x2 & ~x3 & ~x6 & ~x1 & ~x5;
  assign f18 = x4 & x6 & ~x0 & ~x2 & ~x3 & ~x5 & ~x1 & ~x7;
  assign f19 = x0 & x1 & x3 & x5 & ~x2 & ~x14 & ~x15 & ~x13 & ~x12 & ~x11 & ~x10 & ~x9 & ~x8 & ~x6 & ~x7 & ~x4;
  assign f20 = x0 & x4 & x3 & x1 & ~x2 & ~x14 & ~x15 & ~x13 & ~x12 & ~x11 & ~x10 & ~x9 & ~x8 & ~x6 & ~x7 & ~x5;
  assign f21 = ~x11 & ~x12 & ~x3 & ~x2 & ~x0 & x1 & ((x6 & ~x4 & ~x8 & x7 & x5 & (x9 ^ x10) & (x13 ? (~x15 & ~x14) : (~x15 ^ ~x14))) | (~x9 & ~x13 & x4 & x8 & ~x15 & ~x14 & x10 & ~x7 & ~x5));
  assign f22 = ~x11 & ~x12 & ~x3 & ~x2 & ~x0 & x1 & ((x6 & ~x8 & x7 & x4 & x5 & (x9 ^ x10) & (x13 ? (~x15 & ~x14) : (x15 ^ x14))) | (~x13 & ~x15 & x8 & ~x9 & ~x14 & x10 & ~x7 & ~x4 & ~x5));
  assign f23 = ~x3 & ((x0 & ~x1) | (~x2 & ~x0 & x1 & ((~x8 & ~x11 & ~x12 & (x9 ^ x10) & (x13 ? (~x15 & ~x14) : (x15 ^ x14)) & (x6 | ~x5 | (x4 & ~x7))) | (~x5 & x7))));
  assign f24 = x4 & x1 & x3 & x6 & ~x0 & ~x7 & ~x2;
  assign f25 = x4 & x7 & x3 & x1 & ~x0 & ~x6 & ~x2;
  assign f26 = (~x2 & ~x0 & x1 & ((x4 & ((~x5 & x3 & (x6 | x7)) | (~x7 & ~x8 & ~x9 & ~x11 & ~x12 & x10 & ~x3 & (x13 ? (~x15 & ~x14) : (x15 ^ x14))))) | (~x8 & ~x9 & ~x11 & ~x12 & x10 & ~x3 & (x13 ? (~x15 & ~x14) : (x15 ^ x14)) & (x5 ? x6 : ~x7)))) | (~x3 & ~x1 & ~x7 & x0);
  assign f27 = (x7 & ((x4 & x5 & ~x2 & ~x0 & x3 & x1) | (x0 & ~x3 & ~x1))) | (~x2 & ~x0 & x1 & ((~x8 & ~x10 & ~x11 & ~x12 & x9 & ~x3 & (x13 ? (~x15 & ~x14) : (x15 ^ x14)) & ((x6 & x5) | (~x7 & (x4 | ~x5)))) | (x6 & x4 & x5 & x3)));
  assign f28 = ~x3 & ((~x8 & ~x11 & ~x12 & ~x13 & ~x14 & ~x2 & x15 & ~x0 & x1 & ((~x7 & (((x9 | x10) & (x4 | ~x5)) | (x6 & x10))) | (x5 & x6 & (x9 ^ x10)))) | (~x6 & x0 & ~x1));
  assign f29 = ~x8 & ~x11 & ~x12 & ~x15 & ~x14 & ~x3 & ~x2 & ~x0 & x13 & x1 & ((~x7 & (((x9 | x10) & (x4 | ~x5)) | (x6 & x10))) | (x6 & x5 & (x9 ^ x10)));
  assign f30 = ~x3 & ((~x2 & ~x0 & ((~x8 & ~x11 & ~x12 & ~x13 & ~x15 & x14 & x1 & ((~x7 & (((x9 | x10) & (x4 | ~x5)) | (x6 & x10))) | (x6 & x5 & (~x9 ^ ~x10)))) | (x4 & x5 & x7 & ~x1))) | (x6 & x0 & ~x1));
  assign f31 = ~x2 & ~x0 & x1 & ((x4 & x3 & (x6 ? x7 : (x5 & ~x7))) | (~x5 & x7 & ~x3));
  assign f32 = x4 & ((~x3 & ((~x1 & (x0 | (x5 & ~x2 & x7))) | (~x0 & ~x2 & ((~x8 & ~x11 & ~x12 & (x13 ? (~x15 & ~x14) : (x15 ^ x14)) & ((x6 & x5 & x7 & (x9 ^ x10)) | (x1 & ~x7 & (x9 | x10)))) | (~x5 & x1 & x7))))) | (~x6 & x5 & x1 & ~x0 & ~x2 & ~x7 & x3));
  assign f33 = ~x3 & ~x4 & ((x0 & ~x1) | (~x2 & ~x0 & x1 & ((x7 & ~x5) | (~x8 & ~x11 & ~x12 & (x13 ? (~x15 & ~x14) : (x15 ^ x14)) & ((~x5 & (x9 | x10)) | (x6 & (x10 ? (~x7 | ~x9) : x9)))))));
  assign f34 = x4 & x5 & x7 & ~x0 & ~x2 & ~x1 & ~x3;
  assign f35 = ~x1 & ~x3 & ~x2 & ~x0 & x8 & ((x6 & ((x5 & ((x4 & ((x12 & (x13 ? (~x10 & x11) : (x10 & ~x11))) | (x14 & (x15 ? (~x10 & x11) : (x10 & ~x11))))) | (~x10 & ~x11 & ~x4))) | (~x4 & ((~x7 & (x10 ^ x11)) | (~x9 & x7 & ~x5))))) | ((x5 ^ x4) & (~x7 | (~x9 & ~x10 & ~x11))) | (x4 & (x5 ? x7 : ~x6)) | (x7 & ~x6 & ~x5 & (x10 ^ x11)));
  assign f36 = ~x1 & ~x3 & ~x2 & ~x0 & x9 & ((x6 & ((x5 & ((x4 & ((x12 & (x13 ? (~x10 & x11) : (x10 & ~x11))) | (x14 & (x15 ? (~x10 & x11) : (x10 & ~x11))))) | (~x10 & ~x11 & ~x4))) | (~x4 & ((~x7 & (x10 ^ x11)) | (~x8 & x7 & ~x5))))) | ((x5 ^ x4) & (~x7 | (~x8 & ~x10 & ~x11))) | (x4 & (x5 ? x7 : ~x6)) | (x7 & ~x6 & ~x5 & (x10 ^ x11)));
  assign f37 = ~x1 & ~x3 & ~x2 & ~x0 & x10 & ((~x4 & ((~x8 & ((~x9 & ~x11 & ~x6 & x5) | (x9 & x7 & x6 & ~x5))) | (~x7 & (x5 | (~x11 & x6))) | (x8 & ~x9 & x7 & x6 & ~x5))) | (x7 & ((x4 & x5) | (~x11 & ~x6 & ~x5))) | (x4 & ((~x11 & x6 & x5 & ((~x15 & x14) | (~x13 & x12))) | (~x5 & (~x7 | ~x6)))));
  assign f38 = ~x1 & ~x3 & ~x2 & ~x0 & x11 & ((~x4 & ((~x8 & ((~x9 & ~x10 & ~x6 & x5) | (x9 & x7 & x6 & ~x5))) | (~x7 & (x5 | (~x10 & x6))) | (x8 & ~x9 & x7 & x6 & ~x5))) | (x7 & ((x4 & x5) | (~x10 & ~x6 & ~x5))) | (x4 & ((~x5 & (~x7 | ~x6)) | (~x10 & x6 & x5 & ((x15 & x14) | (x12 & x13))))));
  assign f39 = ~x7 & ~x1 & ~x3 & ~x2 & ~x0 & x4 & x6 & x5 & ((x12 & (x13 ? (~x10 & x11) : (x10 & ~x11))) | (x14 & (x15 ? (~x10 & x11) : (x10 & ~x11))));
  assign f40 = ~x7 & ~x11 & ~x12 & ~x3 & ~x2 & ~x0 & x1 & ((~x6 & x4 & x5 & ~x8 & (x9 | x10) & (x13 ? (~x15 & ~x14) : (~x15 ^ ~x14))) | (~x14 & ~x4 & ~x5 & x8 & ~x13 & ~x15 & ~x9 & ~x10));
  assign f41 = x0 & x5 & x7 & x6 & x1 & ~x2 & ~x3 & ~x11 & ~x10 & ~x9 & ~x4 & ~x8;
  assign f42 = ~x1 & ~x5 & ~x4 & ~x3 & ~x2 & ~x0 & (x10 ^ x11) & (x7 ^ x6);
  assign f43 = ~x4 & ~x1 & ~x3 & ~x2 & ~x0 & x6 & ((x7 & ~x5 & (x8 ^ x9)) | (x5 & (~x7 | (~x10 & ~x11))));
  assign f44 = ~x4 & ~x1 & ~x3 & ~x2 & ~x0 & (((x8 ^ x9) & ((~x10 & ~x11 & ~x6 & x5) | (x7 & x6 & ~x5))) | (x5 & (~x7 | (~x6 & ~x8 & ~x9 & (x10 ^ x11)))));
  assign f45 = ~x2 & ~x0 & ((x4 & ((x5 & ((x7 & ~x3 & ~x1) | (x3 & x1 & ~x6 & ~x7))) | (~x8 & ~x11 & ~x12 & x9 & x10 & ~x7 & ~x3 & x1 & (x13 ? (~x15 & ~x14) : (x15 ^ x14))))) | (~x8 & ~x11 & ~x12 & x9 & x10 & ~x7 & ~x3 & x1 & (x6 | ~x5) & (x13 ? (~x15 & ~x14) : (x15 ^ x14))));
endmodule


