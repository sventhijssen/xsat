// Benchmark "top" written by ABC on Fri Mar 31 12:07:43 2023

module top ( 
    pv96_30_, pv96_31_, pv96_10_, pv96_21_, pv138_4_, pv96_11_, pv96_20_,
    pv138_3_, pv138_2_, pv131_18_, pv138_0_, pv131_19_, pv32_7_, pv32_18_,
    pv32_29_, pv64_0_, pv96_9_, pv131_3_, pv131_29_, pv32_6_, pv32_19_,
    pv32_28_, pv64_1_, pv96_8_, pv131_2_, pv131_28_, pv32_5_, pv131_1_,
    pv32_4_, pv131_0_, pv32_3_, pv64_4_, pv96_5_, pv32_2_, pv64_5_,
    pv96_4_, pv32_1_, pv64_2_, pv96_7_, pv32_0_, pv64_3_, pv96_6_,
    pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_, pv97_0_,
    pv131_21_, pv32_11_, pv32_20_, pv64_9_, pv64_18_, pv64_27_, pv96_0_,
    pv131_20_, pv32_12_, pv32_23_, pv32_30_, pv64_6_, pv64_15_, pv64_26_,
    pv96_3_, pv99_0_, pv131_9_, pv131_23_, pv134_0_, pv32_13_, pv32_22_,
    pv32_31_, pv64_7_, pv64_16_, pv64_25_, pv96_2_, pv98_0_, pv131_8_,
    pv131_22_, pv32_14_, pv32_25_, pv131_7_, pv131_25_, pv131_30_,
    pv133_1_, pv32_15_, pv32_24_, pv131_6_, pv131_24_, pv131_31_, pv133_0_,
    pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv131_5_, pv131_27_, pv32_8_,
    pv32_17_, pv32_26_, pv64_29_, pv131_4_, pv131_26_, pv64_20_, pv64_31_,
    pv96_16_, pv96_27_, pv131_16_, pv64_10_, pv96_17_, pv96_26_, pv131_17_,
    pv96_18_, pv96_29_, pv131_14_, pv96_19_, pv96_28_, pv131_15_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv131_12_, pv64_14_, pv64_23_, pv96_13_,
    pv96_22_, pv131_13_, pv64_11_, pv64_22_, pv96_14_, pv96_25_, pv131_10_,
    pv64_12_, pv64_21_, pv64_30_, pv96_15_, pv96_24_, pv131_11_,
    pv198_17_, pv205_3_, pv198_16_, pv205_4_, pv198_19_, pv205_5_,
    pv198_18_, pv205_6_, pv198_8_, pv198_13_, pv198_7_, pv198_12_,
    pv205_0_, pv198_15_, pv205_1_, pv198_9_, pv198_14_, pv205_2_, pv166_7_,
    pv166_10_, pv166_23_, pv198_4_, pv198_22_, pv166_8_, pv166_24_,
    pv198_3_, pv198_23_, pv166_5_, pv166_21_, pv198_6_, pv198_24_,
    pv166_6_, pv166_22_, pv198_5_, pv198_25_, pv166_14_, pv198_0_,
    pv198_26_, pv166_13_, pv166_20_, pv198_27_, pv166_9_, pv166_12_,
    pv198_2_, pv198_28_, pv166_11_, pv198_1_, pv198_29_, pv166_18_,
    pv166_0_, pv166_17_, pv166_16_, pv166_15_, pv166_3_, pv166_27_,
    pv198_31_, pv166_4_, pv198_30_, pv166_1_, pv166_25_, pv198_20_,
    pv166_2_, pv166_19_, pv166_26_, pv198_21_, pv198_11_, pv198_10_  );
  input  pv96_30_, pv96_31_, pv96_10_, pv96_21_, pv138_4_, pv96_11_,
    pv96_20_, pv138_3_, pv138_2_, pv131_18_, pv138_0_, pv131_19_, pv32_7_,
    pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv131_3_, pv131_29_, pv32_6_,
    pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv131_2_, pv131_28_, pv32_5_,
    pv131_1_, pv32_4_, pv131_0_, pv32_3_, pv64_4_, pv96_5_, pv32_2_,
    pv64_5_, pv96_4_, pv32_1_, pv64_2_, pv96_7_, pv32_0_, pv64_3_, pv96_6_,
    pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_, pv97_0_,
    pv131_21_, pv32_11_, pv32_20_, pv64_9_, pv64_18_, pv64_27_, pv96_0_,
    pv131_20_, pv32_12_, pv32_23_, pv32_30_, pv64_6_, pv64_15_, pv64_26_,
    pv96_3_, pv99_0_, pv131_9_, pv131_23_, pv134_0_, pv32_13_, pv32_22_,
    pv32_31_, pv64_7_, pv64_16_, pv64_25_, pv96_2_, pv98_0_, pv131_8_,
    pv131_22_, pv32_14_, pv32_25_, pv131_7_, pv131_25_, pv131_30_,
    pv133_1_, pv32_15_, pv32_24_, pv131_6_, pv131_24_, pv131_31_, pv133_0_,
    pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv131_5_, pv131_27_, pv32_8_,
    pv32_17_, pv32_26_, pv64_29_, pv131_4_, pv131_26_, pv64_20_, pv64_31_,
    pv96_16_, pv96_27_, pv131_16_, pv64_10_, pv96_17_, pv96_26_, pv131_17_,
    pv96_18_, pv96_29_, pv131_14_, pv96_19_, pv96_28_, pv131_15_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv131_12_, pv64_14_, pv64_23_, pv96_13_,
    pv96_22_, pv131_13_, pv64_11_, pv64_22_, pv96_14_, pv96_25_, pv131_10_,
    pv64_12_, pv64_21_, pv64_30_, pv96_15_, pv96_24_, pv131_11_;
  output pv198_17_, pv205_3_, pv198_16_, pv205_4_, pv198_19_, pv205_5_,
    pv198_18_, pv205_6_, pv198_8_, pv198_13_, pv198_7_, pv198_12_,
    pv205_0_, pv198_15_, pv205_1_, pv198_9_, pv198_14_, pv205_2_, pv166_7_,
    pv166_10_, pv166_23_, pv198_4_, pv198_22_, pv166_8_, pv166_24_,
    pv198_3_, pv198_23_, pv166_5_, pv166_21_, pv198_6_, pv198_24_,
    pv166_6_, pv166_22_, pv198_5_, pv198_25_, pv166_14_, pv198_0_,
    pv198_26_, pv166_13_, pv166_20_, pv198_27_, pv166_9_, pv166_12_,
    pv198_2_, pv198_28_, pv166_11_, pv198_1_, pv198_29_, pv166_18_,
    pv166_0_, pv166_17_, pv166_16_, pv166_15_, pv166_3_, pv166_27_,
    pv198_31_, pv166_4_, pv198_30_, pv166_1_, pv166_25_, pv198_20_,
    pv166_2_, pv166_19_, pv166_26_, pv198_21_, pv198_11_, pv198_10_;
  wire new_n_n144_, new_n_n145_, new_n_n196_, new_n_n207_, new_n_n213_,
    new_n_n197_, new_n_n206_, new_n_n148_, new_n_n271_, new_n_n172_,
    new_n_n272_, new_n_n173_, new_n_n250_, new_n_n261_, new_n_n183_,
    new_n_n215_, new_n_n195_, new_n_n157_, new_n_n136_, new_n_n249_,
    new_n_n262_, new_n_n182_, new_n_n216_, new_n_n194_, new_n_n156_,
    new_n_n135_, new_n_n248_, new_n_n155_, new_n_n247_, new_n_n154_,
    new_n_n246_, new_n_n219_, new_n_n191_, new_n_n245_, new_n_n220_,
    new_n_n190_, new_n_n244_, new_n_n217_, new_n_n193_, new_n_n243_,
    new_n_n218_, new_n_n192_, new_n_n253_, new_n_n264_, new_n_n223_,
    new_n_n232_, new_n_n150_, new_n_n187_, new_n_n146_, new_n_n175_,
    new_n_n254_, new_n_n263_, new_n_n224_, new_n_n233_, new_n_n242_,
    new_n_n186_, new_n_n174_, new_n_n255_, new_n_n266_, new_n_n184_,
    new_n_n221_, new_n_n230_, new_n_n241_, new_n_n189_, new_n_n149_,
    new_n_n163_, new_n_n177_, new_n_n141_, new_n_n256_, new_n_n265_,
    new_n_n185_, new_n_n222_, new_n_n231_, new_n_n240_, new_n_n188_,
    new_n_n147_, new_n_n162_, new_n_n176_, new_n_n257_, new_n_n268_,
    new_n_n161_, new_n_n179_, new_n_n137_, new_n_n140_, new_n_n258_,
    new_n_n267_, new_n_n160_, new_n_n178_, new_n_n138_, new_n_n139_,
    new_n_n252_, new_n_n259_, new_n_n270_, new_n_n234_, new_n_n159_,
    new_n_n181_, new_n_n251_, new_n_n260_, new_n_n269_, new_n_n151_,
    new_n_n158_, new_n_n180_, new_n_n235_, new_n_n153_, new_n_n202_,
    new_n_n214_, new_n_n170_, new_n_n225_, new_n_n203_, new_n_n212_,
    new_n_n171_, new_n_n204_, new_n_n143_, new_n_n168_, new_n_n205_,
    new_n_n142_, new_n_n169_, new_n_n228_, new_n_n239_, new_n_n198_,
    new_n_n209_, new_n_n166_, new_n_n229_, new_n_n238_, new_n_n199_,
    new_n_n208_, new_n_n167_, new_n_n226_, new_n_n237_, new_n_n200_,
    new_n_n211_, new_n_n164_, new_n_n227_, new_n_n236_, new_n_n152_,
    new_n_n201_, new_n_n210_, new_n_n165_, new_nv212_, new_nv223_,
    new_nv234_, new_n_n130_, new_nv257_, new_n_n108_, new_nv300_,
    new_nv311_, new_nv324_, new_nv335_, new_nv346_, new_nv372_, new_n_n83_,
    new_nv383_, new_nv423_, new_nv434_, new_nv445_, new_nv213_, new_nv222_,
    new_nv235_, new_nv240_, new_nv252_, new_nv263_, new_nv299_, new_nv312_,
    new_nv323_, new_nv336_, new_nv345_, new_n_n88_, new_nv377_, new_n_n77_,
    new_nv422_, new_nv435_, new_nv444_, new_nv214_, new_nv225_, new_nv232_,
    new_n_n131_, new_n_n118_, new_nv258_, new_nv298_, new_nv313_,
    new_nv326_, new_nv333_, new_nv344_, new_nv362_, new_n_n93_, new_nv384_,
    new_nv425_, new_nv432_, new_nv443_, new_nv215_, new_nv224_, new_nv233_,
    new_nv239_, new_nv253_, new_n_n113_, new_nv262_, new_nv314_,
    new_nv325_, new_nv334_, new_nv343_, new_n_n98_, new_nv367_, new_n_n76_,
    new_nv424_, new_nv433_, new_nv442_, new_nv216_, new_nv227_,
    new_n_n128_, new_nv248_, new_nv315_, new_nv328_, new_nv339_,
    new_nv350_, new_n_n103_, new_nv385_, new_nv427_, new_nv438_,
    new_nv449_, new_n_n7_, new_nv217_, new_nv226_, new_nv243_, new_n_n123_,
    new_nv316_, new_nv327_, new_nv349_, new_nv351_, new_nv357_, new_n_n75_,
    new_nv426_, new_nv439_, new_nv448_, new_nv236_, new_n_n129_,
    new_nv247_, new_nv317_, new_nv337_, new_nv348_, new_nv418_, new_nv429_,
    new_nv436_, new_nv447_, new_n_n134_, new_nv241_, new_nv242_,
    new_nv329_, new_nv338_, new_nv347_, new_nv419_, new_nv428_, new_nv437_,
    new_nv446_, new_n_n126_, new_nv250_, new_n_n115_, new_nv261_,
    new_nv297_, new_nv354_, new_n_n101_, new_nv365_, new_n_n90_,
    new_nv376_, new_n_n79_, new_n_n3_, new_nv245_, new_n_n121_, new_nv256_,
    new_n_n110_, new_nv307_, new_n_n106_, new_nv359_, new_n_n95_,
    new_nv370_, new_n_n84_, new_nv381_, new_n_n4_, new_n_n127_, new_nv249_,
    new_n_n114_, new_nv295_, new_nv306_, new_nv352_, new_n_n102_,
    new_nv366_, new_n_n89_, new_nv375_, new_n_n80_, new_n_n5_, new_nv244_,
    new_n_n122_, new_n_n109_, new_nv296_, new_nv305_, new_nv353_,
    new_nv358_, new_n_n94_, new_nv371_, new_n_n85_, new_nv380_, new_n_n6_,
    new_nv208_, new_nv219_, new_nv230_, new_n_n132_, new_n_n124_,
    new_n_n117_, new_nv259_, new_nv293_, new_nv304_, new_nv318_,
    new_nv331_, new_nv342_, new_nv356_, new_n_n99_, new_nv363_, new_n_n92_,
    new_nv374_, new_n_n81_, new_nv430_, new_nv441_, new_nv452_, new_nv209_,
    new_nv218_, new_nv231_, new_nv238_, new_n_n119_, new_nv254_,
    new_n_n112_, new_nv294_, new_nv303_, new_nv308_, new_nv332_,
    new_nv341_, new_n_n104_, new_nv361_, new_n_n97_, new_nv368_,
    new_n_n86_, new_nv379_, new_nv431_, new_nv440_, new_nv453_, new_nv210_,
    new_nv221_, new_nv228_, new_n_n133_, new_n_n125_, new_nv251_,
    new_n_n116_, new_nv260_, new_n_n107_, new_nv302_, new_nv309_,
    new_nv322_, new_nv340_, new_nv355_, new_n_n100_, new_nv364_,
    new_n_n91_, new_nv373_, new_n_n82_, new_nv382_, new_nv421_, new_nv481_,
    new_nv211_, new_nv220_, new_nv229_, new_nv237_, new_nv246_,
    new_n_n120_, new_nv255_, new_n_n111_, new_nv292_, new_nv301_,
    new_nv310_, new_nv319_, new_nv330_, new_n_n105_, new_nv360_,
    new_n_n96_, new_nv369_, new_n_n87_, new_nv378_, new_n_n78_, new_nv420_,
    new_n_n2_, new_nv458_, new_nv465_, new_nv479_, new_n_n59_, new_n_n48_,
    new_nv457_, new_n_n70_, new_nv478_, new_n_n58_, new_n_n49_, new_nv456_,
    new_nv466_, new_nv482_, new_n_n61_, new_n_n50_, new_nv455_, new_n_n69_,
    new_nv480_, new_n_n60_, new_n_n51_, new_nv450_, new_nv454_, new_n_n41_,
    new_n_n30_, new_n_n19_, new_n_n8_, new_nv451_, new_n_n40_, new_n_n31_,
    new_n_n18_, new_n_n9_, new_n_n39_, new_n_n28_, new_n_n21_, new_n_n10_,
    new_n_n38_, new_n_n29_, new_n_n20_, new_n_n11_, new_n_n67_, new_n_n56_,
    new_n_n45_, new_n_n34_, new_n_n23_, new_n_n12_, new_n_n66_, new_n_n57_,
    new_n_n44_, new_n_n35_, new_n_n22_, new_n_n13_, new_nv462_, new_n_n68_,
    new_n_n43_, new_n_n32_, new_n_n25_, new_n_n14_, new_n_n73_, new_nv467_,
    new_n_n42_, new_n_n33_, new_n_n24_, new_n_n15_, new_n_n74_, new_nv463_,
    new_nv475_, new_n_n63_, new_n_n52_, new_n_n27_, new_n_n16_, new_nv461_,
    new_n_n72_, new_nv474_, new_n_n62_, new_n_n53_, new_n_n26_, new_n_n17_,
    new_nv460_, new_nv464_, new_nv477_, new_n_n65_, new_n_n54_, new_n_n47_,
    new_n_n36_, new_nv459_, new_n_n71_, new_nv476_, new_n_n64_, new_n_n55_,
    new_n_n46_, new_n_n37_;
  assign new_n_n144_ = pv96_30_;
  assign pv198_17_ = new_n_n92_;
  assign pv205_3_ = new_n_n71_;
  assign new_n_n145_ = pv96_31_;
  assign pv198_16_ = new_n_n91_;
  assign pv205_4_ = new_n_n72_;
  assign new_n_n196_ = pv96_10_;
  assign new_n_n207_ = pv96_21_;
  assign new_n_n213_ = pv138_4_;
  assign pv198_19_ = new_n_n94_;
  assign pv205_5_ = new_n_n73_;
  assign new_n_n197_ = pv96_11_;
  assign new_n_n206_ = pv96_20_;
  assign new_n_n148_ = pv138_3_;
  assign pv198_18_ = new_n_n93_;
  assign pv205_6_ = new_n_n74_;
  assign new_n_n271_ = pv138_2_;
  assign pv198_8_ = new_n_n83_;
  assign pv198_13_ = new_n_n88_;
  assign pv198_7_ = new_n_n82_;
  assign pv198_12_ = new_n_n87_;
  assign pv205_0_ = new_n_n68_;
  assign new_n_n172_ = pv131_18_;
  assign new_n_n272_ = pv138_0_;
  assign pv198_15_ = new_n_n90_;
  assign pv205_1_ = new_n_n69_;
  assign new_n_n173_ = pv131_19_;
  assign pv198_9_ = new_n_n84_;
  assign pv198_14_ = new_n_n89_;
  assign pv205_2_ = new_n_n70_;
  assign new_n_n250_ = pv32_7_;
  assign new_n_n261_ = pv32_18_;
  assign new_n_n183_ = pv32_29_;
  assign new_n_n215_ = pv64_0_;
  assign new_n_n195_ = pv96_9_;
  assign new_n_n157_ = pv131_3_;
  assign new_n_n136_ = pv131_29_;
  assign pv166_7_ = new_n_n114_;
  assign pv166_10_ = new_n_n117_;
  assign pv166_23_ = new_n_n130_;
  assign pv198_4_ = new_n_n79_;
  assign pv198_22_ = new_n_n97_;
  assign new_n_n249_ = pv32_6_;
  assign new_n_n262_ = pv32_19_;
  assign new_n_n182_ = pv32_28_;
  assign new_n_n216_ = pv64_1_;
  assign new_n_n194_ = pv96_8_;
  assign new_n_n156_ = pv131_2_;
  assign new_n_n135_ = pv131_28_;
  assign pv166_8_ = new_n_n115_;
  assign pv166_24_ = new_n_n131_;
  assign pv198_3_ = new_n_n78_;
  assign pv198_23_ = new_n_n98_;
  assign new_n_n248_ = pv32_5_;
  assign new_n_n155_ = pv131_1_;
  assign pv166_5_ = new_n_n112_;
  assign pv166_21_ = new_n_n128_;
  assign pv198_6_ = new_n_n81_;
  assign pv198_24_ = new_n_n99_;
  assign new_n_n247_ = pv32_4_;
  assign new_n_n154_ = pv131_0_;
  assign pv166_6_ = new_n_n113_;
  assign pv166_22_ = new_n_n129_;
  assign pv198_5_ = new_n_n80_;
  assign pv198_25_ = new_n_n100_;
  assign new_n_n246_ = pv32_3_;
  assign new_n_n219_ = pv64_4_;
  assign new_n_n191_ = pv96_5_;
  assign pv166_14_ = new_n_n121_;
  assign pv198_0_ = new_n_n75_;
  assign pv198_26_ = new_n_n101_;
  assign new_n_n245_ = pv32_2_;
  assign new_n_n220_ = pv64_5_;
  assign new_n_n190_ = pv96_4_;
  assign pv166_13_ = new_n_n120_;
  assign pv166_20_ = new_n_n127_;
  assign pv198_27_ = new_n_n102_;
  assign new_n_n244_ = pv32_1_;
  assign new_n_n217_ = pv64_2_;
  assign new_n_n193_ = pv96_7_;
  assign pv166_9_ = new_n_n116_;
  assign pv166_12_ = new_n_n119_;
  assign pv198_2_ = new_n_n77_;
  assign pv198_28_ = new_n_n103_;
  assign new_n_n243_ = pv32_0_;
  assign new_n_n218_ = pv64_3_;
  assign new_n_n192_ = pv96_6_;
  assign pv166_11_ = new_n_n118_;
  assign pv198_1_ = new_n_n76_;
  assign pv198_29_ = new_n_n104_;
  assign new_n_n253_ = pv32_10_;
  assign new_n_n264_ = pv32_21_;
  assign new_n_n223_ = pv64_8_;
  assign new_n_n232_ = pv64_17_;
  assign new_n_n150_ = pv64_28_;
  assign new_n_n187_ = pv96_1_;
  assign new_n_n146_ = pv97_0_;
  assign new_n_n175_ = pv131_21_;
  assign pv166_18_ = new_n_n125_;
  assign new_n_n254_ = pv32_11_;
  assign new_n_n263_ = pv32_20_;
  assign new_n_n224_ = pv64_9_;
  assign new_n_n233_ = pv64_18_;
  assign new_n_n242_ = pv64_27_;
  assign new_n_n186_ = pv96_0_;
  assign new_n_n174_ = pv131_20_;
  assign pv166_0_ = new_n_n107_;
  assign pv166_17_ = new_n_n124_;
  assign new_n_n255_ = pv32_12_;
  assign new_n_n266_ = pv32_23_;
  assign new_n_n184_ = pv32_30_;
  assign new_n_n221_ = pv64_6_;
  assign new_n_n230_ = pv64_15_;
  assign new_n_n241_ = pv64_26_;
  assign new_n_n189_ = pv96_3_;
  assign new_n_n149_ = pv99_0_;
  assign new_n_n163_ = pv131_9_;
  assign new_n_n177_ = pv131_23_;
  assign new_n_n141_ = pv134_0_;
  assign pv166_16_ = new_n_n123_;
  assign new_n_n256_ = pv32_13_;
  assign new_n_n265_ = pv32_22_;
  assign new_n_n185_ = pv32_31_;
  assign new_n_n222_ = pv64_7_;
  assign new_n_n231_ = pv64_16_;
  assign new_n_n240_ = pv64_25_;
  assign new_n_n188_ = pv96_2_;
  assign new_n_n147_ = pv98_0_;
  assign new_n_n162_ = pv131_8_;
  assign new_n_n176_ = pv131_22_;
  assign pv166_15_ = new_n_n122_;
  assign new_n_n257_ = pv32_14_;
  assign new_n_n268_ = pv32_25_;
  assign new_n_n161_ = pv131_7_;
  assign new_n_n179_ = pv131_25_;
  assign new_n_n137_ = pv131_30_;
  assign new_n_n140_ = pv133_1_;
  assign pv166_3_ = new_n_n110_;
  assign pv166_27_ = new_n_n134_;
  assign pv198_31_ = new_n_n106_;
  assign new_n_n258_ = pv32_15_;
  assign new_n_n267_ = pv32_24_;
  assign new_n_n160_ = pv131_6_;
  assign new_n_n178_ = pv131_24_;
  assign new_n_n138_ = pv131_31_;
  assign new_n_n139_ = pv133_0_;
  assign pv166_4_ = new_n_n111_;
  assign pv198_30_ = new_n_n105_;
  assign new_n_n252_ = pv32_9_;
  assign new_n_n259_ = pv32_16_;
  assign new_n_n270_ = pv32_27_;
  assign new_n_n234_ = pv64_19_;
  assign new_n_n159_ = pv131_5_;
  assign new_n_n181_ = pv131_27_;
  assign pv166_1_ = new_n_n108_;
  assign pv166_25_ = new_n_n132_;
  assign pv198_20_ = new_n_n95_;
  assign new_n_n251_ = pv32_8_;
  assign new_n_n260_ = pv32_17_;
  assign new_n_n269_ = pv32_26_;
  assign new_n_n151_ = pv64_29_;
  assign new_n_n158_ = pv131_4_;
  assign new_n_n180_ = pv131_26_;
  assign pv166_2_ = new_n_n109_;
  assign pv166_19_ = new_n_n126_;
  assign pv166_26_ = new_n_n133_;
  assign pv198_21_ = new_n_n96_;
  assign new_n_n235_ = pv64_20_;
  assign new_n_n153_ = pv64_31_;
  assign new_n_n202_ = pv96_16_;
  assign new_n_n214_ = pv96_27_;
  assign new_n_n170_ = pv131_16_;
  assign new_n_n225_ = pv64_10_;
  assign new_n_n203_ = pv96_17_;
  assign new_n_n212_ = pv96_26_;
  assign new_n_n171_ = pv131_17_;
  assign new_n_n204_ = pv96_18_;
  assign new_n_n143_ = pv96_29_;
  assign new_n_n168_ = pv131_14_;
  assign pv198_11_ = new_n_n86_;
  assign new_n_n205_ = pv96_19_;
  assign new_n_n142_ = pv96_28_;
  assign new_n_n169_ = pv131_15_;
  assign pv198_10_ = new_n_n85_;
  assign new_n_n228_ = pv64_13_;
  assign new_n_n239_ = pv64_24_;
  assign new_n_n198_ = pv96_12_;
  assign new_n_n209_ = pv96_23_;
  assign new_n_n166_ = pv131_12_;
  assign new_n_n229_ = pv64_14_;
  assign new_n_n238_ = pv64_23_;
  assign new_n_n199_ = pv96_13_;
  assign new_n_n208_ = pv96_22_;
  assign new_n_n167_ = pv131_13_;
  assign new_n_n226_ = pv64_11_;
  assign new_n_n237_ = pv64_22_;
  assign new_n_n200_ = pv96_14_;
  assign new_n_n211_ = pv96_25_;
  assign new_n_n164_ = pv131_10_;
  assign new_n_n227_ = pv64_12_;
  assign new_n_n236_ = pv64_21_;
  assign new_n_n152_ = pv64_30_;
  assign new_n_n201_ = pv96_15_;
  assign new_n_n210_ = pv96_24_;
  assign new_n_n165_ = pv131_11_;
  assign new_nv212_ = new_n_n266_ & new_nv453_ & new_nv452_;
  assign new_nv223_ = new_n_n255_ & new_nv453_ & new_nv452_;
  assign new_nv234_ = new_n_n244_ & new_nv453_ & new_nv452_;
  assign new_n_n130_ = new_nv296_ | new_nv240_ | new_nv212_;
  assign new_nv257_ = new_n_n221_ & new_nv453_ & new_n_n272_;
  assign new_n_n108_ = new_nv318_ | new_nv262_ | new_nv234_;
  assign new_nv300_ = new_n_n21_ & new_n_n271_ & new_n_n272_;
  assign new_nv311_ = new_n_n10_ & new_n_n271_ & new_n_n272_;
  assign new_nv324_ = new_n_n211_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv335_ = new_n_n200_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv346_ = new_n_n189_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv372_ = new_n_n163_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n83_ = new_nv345_ | new_nv441_ | new_nv377_ | new_nv451_;
  assign new_nv383_ = new_n_n152_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_nv423_ = new_n_n56_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv434_ = new_n_n45_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv445_ = new_n_n34_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv213_ = new_n_n265_ & new_nv453_ & new_nv452_;
  assign new_nv222_ = new_n_n256_ & new_nv453_ & new_nv452_;
  assign new_nv235_ = new_n_n243_ & new_nv453_ & new_nv452_;
  assign new_nv240_ = new_n_n238_ & new_nv453_ & new_n_n272_;
  assign new_nv252_ = new_n_n226_ & new_nv453_ & new_n_n272_;
  assign new_nv263_ = new_n_n215_ & new_nv453_ & new_n_n272_;
  assign new_nv299_ = new_n_n22_ & new_n_n271_ & new_n_n272_;
  assign new_nv312_ = new_n_n9_ & new_n_n271_ & new_n_n272_;
  assign new_nv323_ = new_n_n212_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv336_ = new_n_n199_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv345_ = new_n_n190_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_n_n88_ = new_nv340_ | new_nv436_ | new_nv372_ | new_nv451_;
  assign new_nv377_ = new_n_n158_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n77_ = new_nv351_ | new_nv447_ | new_nv383_ | new_nv451_;
  assign new_nv422_ = new_n_n57_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv435_ = new_n_n44_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv444_ = new_n_n35_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv214_ = new_n_n264_ & new_nv453_ & new_nv452_;
  assign new_nv225_ = new_n_n253_ & new_nv453_ & new_nv452_;
  assign new_nv232_ = new_n_n246_ & new_nv453_ & new_nv452_;
  assign new_n_n131_ = new_nv295_ | new_nv239_ | new_nv211_;
  assign new_n_n118_ = new_nv308_ | new_nv252_ | new_nv224_;
  assign new_nv258_ = new_n_n220_ & new_nv453_ & new_n_n272_;
  assign new_nv298_ = new_n_n23_ & new_n_n271_ & new_n_n272_;
  assign new_nv313_ = new_n_n8_ & new_n_n271_ & new_n_n272_;
  assign new_nv326_ = new_n_n209_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv333_ = new_n_n202_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv344_ = new_n_n191_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv362_ = new_n_n173_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n93_ = new_nv335_ | new_nv431_ | new_nv367_ | new_nv451_;
  assign new_nv384_ = new_n_n151_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_nv425_ = new_n_n54_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv432_ = new_n_n47_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv443_ = new_n_n36_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv215_ = new_n_n263_ & new_nv453_ & new_nv452_;
  assign new_nv224_ = new_n_n254_ & new_nv453_ & new_nv452_;
  assign new_nv233_ = new_n_n245_ & new_nv453_ & new_nv452_;
  assign new_nv239_ = new_n_n239_ & new_nv453_ & new_n_n272_;
  assign new_nv253_ = new_n_n225_ & new_nv453_ & new_n_n272_;
  assign new_n_n113_ = new_nv313_ | new_nv257_ | new_nv229_;
  assign new_nv262_ = new_n_n216_ & new_nv453_ & new_n_n272_;
  assign new_nv314_ = new_n_n7_ & new_n_n271_ & new_n_n272_;
  assign new_nv325_ = new_n_n210_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv334_ = new_n_n201_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv343_ = new_n_n192_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_n_n98_ = new_nv330_ | new_nv426_ | new_nv362_ | new_nv451_;
  assign new_nv367_ = new_n_n168_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n76_ = new_nv352_ | new_nv448_ | new_nv384_ | new_nv451_;
  assign new_nv424_ = new_n_n55_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv433_ = new_n_n46_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv442_ = new_n_n37_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv216_ = new_n_n262_ & new_nv453_ & new_nv452_;
  assign new_nv227_ = new_n_n251_ & new_nv453_ & new_nv452_;
  assign new_n_n128_ = new_nv298_ | new_nv242_ | new_nv214_;
  assign new_nv248_ = new_n_n230_ & new_nv453_ & new_n_n272_;
  assign new_nv315_ = new_n_n6_ & new_n_n271_ & new_n_n272_;
  assign new_nv328_ = new_n_n207_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv339_ = new_n_n196_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv350_ = new_n_n185_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_n_n103_ = new_nv325_ | new_nv421_ | new_nv357_ | new_nv451_;
  assign new_nv385_ = new_n_n150_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_nv427_ = new_n_n52_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv438_ = new_n_n41_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv449_ = new_n_n30_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_n_n7_ = ~new_n_n220_;
  assign new_nv217_ = new_n_n261_ & new_nv453_ & new_nv452_;
  assign new_nv226_ = new_n_n252_ & new_nv453_ & new_nv452_;
  assign new_nv243_ = new_n_n235_ & new_nv453_ & new_n_n272_;
  assign new_n_n123_ = new_nv303_ | new_nv247_ | new_nv219_;
  assign new_nv316_ = new_n_n5_ & new_n_n271_ & new_n_n272_;
  assign new_nv327_ = new_n_n208_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv349_ = new_n_n186_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv351_ = new_n_n184_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv357_ = new_n_n178_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n75_ = new_nv353_ | new_nv449_ | new_nv385_ | new_nv451_;
  assign new_nv426_ = new_n_n53_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv439_ = new_n_n40_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv448_ = new_n_n31_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv236_ = new_n_n242_ & new_nv453_ & new_n_n272_;
  assign new_n_n129_ = new_nv297_ | new_nv241_ | new_nv213_;
  assign new_nv247_ = new_n_n231_ & new_nv453_ & new_n_n272_;
  assign new_nv317_ = new_n_n4_ & new_n_n271_ & new_n_n272_;
  assign new_nv337_ = new_n_n198_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv348_ = new_n_n187_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv418_ = new_n_n61_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv429_ = new_n_n50_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv436_ = new_n_n43_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv447_ = new_n_n32_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_n_n134_ = new_nv292_ | new_nv236_ | new_nv208_;
  assign new_nv241_ = new_n_n237_ & new_nv453_ & new_n_n272_;
  assign new_nv242_ = new_n_n236_ & new_nv453_ & new_n_n272_;
  assign new_nv329_ = new_n_n206_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv338_ = new_n_n197_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv347_ = new_n_n188_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv419_ = new_n_n60_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv428_ = new_n_n51_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv437_ = new_n_n42_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv446_ = new_n_n33_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_n_n126_ = new_nv300_ | new_nv244_ | new_nv216_;
  assign new_nv250_ = new_n_n228_ & new_nv453_ & new_n_n272_;
  assign new_n_n115_ = new_nv311_ | new_nv255_ | new_nv227_;
  assign new_nv261_ = new_n_n217_ & new_nv453_ & new_n_n272_;
  assign new_nv297_ = new_n_n24_ & new_n_n271_ & new_n_n272_;
  assign new_nv354_ = new_n_n181_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n101_ = new_nv327_ | new_nv423_ | new_nv359_ | new_nv451_;
  assign new_nv365_ = new_n_n170_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n90_ = new_nv338_ | new_nv434_ | new_nv370_ | new_nv451_;
  assign new_nv376_ = new_n_n159_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n79_ = new_nv349_ | new_nv445_ | new_nv381_ | new_nv451_;
  assign new_n_n3_ = ~new_n_n216_;
  assign new_nv245_ = new_n_n233_ & new_nv453_ & new_n_n272_;
  assign new_n_n121_ = new_nv305_ | new_nv249_ | new_nv221_;
  assign new_nv256_ = new_n_n222_ & new_nv453_ & new_n_n272_;
  assign new_n_n110_ = new_nv316_ | new_nv260_ | new_nv232_;
  assign new_nv307_ = new_n_n14_ & new_n_n271_ & new_n_n272_;
  assign new_n_n106_ = new_nv322_ | new_nv418_ | new_nv354_ | new_nv451_;
  assign new_nv359_ = new_n_n176_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n95_ = new_nv333_ | new_nv429_ | new_nv365_ | new_nv451_;
  assign new_nv370_ = new_n_n165_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n84_ = new_nv344_ | new_nv440_ | new_nv376_ | new_nv451_;
  assign new_nv381_ = new_n_n154_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n4_ = ~new_n_n217_;
  assign new_n_n127_ = new_nv299_ | new_nv243_ | new_nv215_;
  assign new_nv249_ = new_n_n229_ & new_nv453_ & new_n_n272_;
  assign new_n_n114_ = new_nv312_ | new_nv256_ | new_nv228_;
  assign new_nv295_ = new_n_n26_ & new_n_n271_ & new_n_n272_;
  assign new_nv306_ = new_n_n15_ & new_n_n271_ & new_n_n272_;
  assign new_nv352_ = new_n_n183_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_n_n102_ = new_nv326_ | new_nv422_ | new_nv358_ | new_nv451_;
  assign new_nv366_ = new_n_n169_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n89_ = new_nv339_ | new_nv435_ | new_nv371_ | new_nv451_;
  assign new_nv375_ = new_n_n160_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n80_ = new_nv348_ | new_nv444_ | new_nv380_ | new_nv451_;
  assign new_n_n5_ = ~new_n_n218_;
  assign new_nv244_ = new_n_n234_ & new_nv453_ & new_n_n272_;
  assign new_n_n122_ = new_nv304_ | new_nv248_ | new_nv220_;
  assign new_n_n109_ = new_nv317_ | new_nv261_ | new_nv233_;
  assign new_nv296_ = new_n_n25_ & new_n_n271_ & new_n_n272_;
  assign new_nv305_ = new_n_n16_ & new_n_n271_ & new_n_n272_;
  assign new_nv353_ = new_n_n182_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv358_ = new_n_n177_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n94_ = new_nv334_ | new_nv430_ | new_nv366_ | new_nv451_;
  assign new_nv371_ = new_n_n164_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n85_ = new_nv343_ | new_nv439_ | new_nv375_ | new_nv451_;
  assign new_nv380_ = new_n_n155_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n6_ = ~new_n_n219_;
  assign new_nv208_ = new_n_n270_ & new_nv453_ & new_nv452_;
  assign new_nv219_ = new_n_n259_ & new_nv453_ & new_nv452_;
  assign new_nv230_ = new_n_n248_ & new_nv453_ & new_nv452_;
  assign new_n_n132_ = new_nv294_ | new_nv238_ | new_nv210_;
  assign new_n_n124_ = new_nv302_ | new_nv246_ | new_nv218_;
  assign new_n_n117_ = new_nv309_ | new_nv253_ | new_nv225_;
  assign new_nv259_ = new_n_n219_ & new_nv453_ & new_n_n272_;
  assign new_nv293_ = new_n_n28_ & new_n_n271_ & new_n_n272_;
  assign new_nv304_ = new_n_n17_ & new_n_n271_ & new_n_n272_;
  assign new_nv318_ = new_n_n3_ & new_n_n271_ & new_n_n272_;
  assign new_nv331_ = new_n_n204_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv342_ = new_n_n193_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv356_ = new_n_n179_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n99_ = new_nv329_ | new_nv425_ | new_nv361_ | new_nv451_;
  assign new_nv363_ = new_n_n172_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n92_ = new_nv336_ | new_nv432_ | new_nv368_ | new_nv451_;
  assign new_nv374_ = new_n_n161_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n81_ = new_nv347_ | new_nv443_ | new_nv379_ | new_nv451_;
  assign new_nv430_ = new_n_n49_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv441_ = new_n_n38_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv452_ = ~new_n_n272_;
  assign new_nv209_ = new_n_n269_ & new_nv453_ & new_nv452_;
  assign new_nv218_ = new_n_n260_ & new_nv453_ & new_nv452_;
  assign new_nv231_ = new_n_n247_ & new_nv453_ & new_nv452_;
  assign new_nv238_ = new_n_n240_ & new_nv453_ & new_n_n272_;
  assign new_n_n119_ = new_nv307_ | new_nv251_ | new_nv223_;
  assign new_nv254_ = new_n_n224_ & new_nv453_ & new_n_n272_;
  assign new_n_n112_ = new_nv314_ | new_nv258_ | new_nv230_;
  assign new_nv294_ = new_n_n27_ & new_n_n271_ & new_n_n272_;
  assign new_nv303_ = new_n_n18_ & new_n_n271_ & new_n_n272_;
  assign new_nv308_ = new_n_n13_ & new_n_n271_ & new_n_n272_;
  assign new_nv332_ = new_n_n203_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv341_ = new_n_n194_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_n_n104_ = new_nv324_ | new_nv420_ | new_nv356_ | new_nv451_;
  assign new_nv361_ = new_n_n174_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n97_ = new_nv331_ | new_nv427_ | new_nv363_ | new_nv451_;
  assign new_nv368_ = new_n_n167_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n86_ = new_nv342_ | new_nv438_ | new_nv374_ | new_nv451_;
  assign new_nv379_ = new_n_n156_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_nv431_ = new_n_n48_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv440_ = new_n_n39_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv453_ = ~new_n_n271_;
  assign new_nv210_ = new_n_n268_ & new_nv453_ & new_nv452_;
  assign new_nv221_ = new_n_n257_ & new_nv453_ & new_nv452_;
  assign new_nv228_ = new_n_n250_ & new_nv453_ & new_nv452_;
  assign new_n_n133_ = new_nv293_ | new_nv237_ | new_nv209_;
  assign new_n_n125_ = new_nv301_ | new_nv245_ | new_nv217_;
  assign new_nv251_ = new_n_n227_ & new_nv453_ & new_n_n272_;
  assign new_n_n116_ = new_nv310_ | new_nv254_ | new_nv226_;
  assign new_nv260_ = new_n_n218_ & new_nv453_ & new_n_n272_;
  assign new_n_n107_ = new_nv319_ | new_nv263_ | new_nv235_;
  assign new_nv302_ = new_n_n19_ & new_n_n271_ & new_n_n272_;
  assign new_nv309_ = new_n_n12_ & new_n_n271_ & new_n_n272_;
  assign new_nv322_ = new_n_n214_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv340_ = new_n_n195_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_nv355_ = new_n_n180_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n100_ = new_nv328_ | new_nv424_ | new_nv360_ | new_nv451_;
  assign new_nv364_ = new_n_n171_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n91_ = new_nv337_ | new_nv433_ | new_nv369_ | new_nv451_;
  assign new_nv373_ = new_n_n162_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n82_ = new_nv346_ | new_nv442_ | new_nv378_ | new_nv451_;
  assign new_nv382_ = new_n_n153_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_nv421_ = new_n_n58_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_nv481_ = ~new_n_n148_;
  assign new_nv211_ = new_n_n267_ & new_nv453_ & new_nv452_;
  assign new_nv220_ = new_n_n258_ & new_nv453_ & new_nv452_;
  assign new_nv229_ = new_n_n249_ & new_nv453_ & new_nv452_;
  assign new_nv237_ = new_n_n241_ & new_nv453_ & new_n_n272_;
  assign new_nv246_ = new_n_n232_ & new_nv453_ & new_n_n272_;
  assign new_n_n120_ = new_nv306_ | new_nv250_ | new_nv222_;
  assign new_nv255_ = new_n_n223_ & new_nv453_ & new_n_n272_;
  assign new_n_n111_ = new_nv315_ | new_nv259_ | new_nv231_;
  assign new_nv292_ = new_n_n29_ & new_n_n271_ & new_n_n272_;
  assign new_nv301_ = new_n_n20_ & new_n_n271_ & new_n_n272_;
  assign new_nv310_ = new_n_n11_ & new_n_n271_ & new_n_n272_;
  assign new_nv319_ = new_n_n2_ & new_n_n271_ & new_n_n272_;
  assign new_nv330_ = new_n_n205_ & new_nv453_ & new_n_n213_ & new_nv452_;
  assign new_n_n105_ = new_nv323_ | new_nv419_ | new_nv355_ | new_nv451_;
  assign new_nv360_ = new_n_n175_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n96_ = new_nv332_ | new_nv428_ | new_nv364_ | new_nv451_;
  assign new_nv369_ = new_n_n166_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n87_ = new_nv341_ | new_nv437_ | new_nv373_ | new_nv451_;
  assign new_nv378_ = new_n_n157_ & new_nv453_ & new_n_n213_ & new_n_n272_;
  assign new_n_n78_ = new_nv350_ | new_nv446_ | new_nv382_ | new_nv451_;
  assign new_nv420_ = new_n_n59_ & new_n_n271_ & new_n_n213_ & new_n_n272_;
  assign new_n_n2_ = ~new_n_n215_;
  assign new_nv458_ = new_n_n144_ & new_nv453_ & new_n_n148_ & new_nv452_;
  assign new_nv465_ = new_n_n137_ & new_nv453_ & new_n_n148_ & new_n_n272_;
  assign new_nv479_ = new_n_n63_ & new_n_n271_ & new_n_n148_ & new_n_n272_;
  assign new_n_n59_ = ~new_n_n179_;
  assign new_n_n48_ = ~new_n_n168_;
  assign new_nv457_ = new_n_n145_ & new_nv453_ & new_n_n148_ & new_nv452_;
  assign new_n_n70_ = new_nv458_ | new_nv478_ | new_nv465_ | new_nv482_;
  assign new_nv478_ = new_n_n64_ & new_n_n271_ & new_n_n148_ & new_n_n272_;
  assign new_n_n58_ = ~new_n_n178_;
  assign new_n_n49_ = ~new_n_n169_;
  assign new_nv456_ = new_n_n146_ & new_nv453_ & new_n_n148_ & new_nv452_;
  assign new_nv466_ = new_n_n136_ & new_nv453_ & new_n_n148_ & new_n_n272_;
  assign new_nv482_ = new_nv481_ & new_n_n271_;
  assign new_n_n61_ = ~new_n_n181_;
  assign new_n_n50_ = ~new_n_n170_;
  assign new_nv455_ = new_n_n147_ & new_nv453_ & new_n_n148_ & new_nv452_;
  assign new_n_n69_ = new_nv459_ | new_nv479_ | new_nv466_ | new_nv482_;
  assign new_nv480_ = new_n_n62_ & new_n_n271_ & new_n_n148_ & new_n_n272_;
  assign new_n_n60_ = ~new_n_n180_;
  assign new_n_n51_ = ~new_n_n171_;
  assign new_nv450_ = ~new_n_n213_;
  assign new_nv454_ = new_n_n149_ & new_nv453_ & new_n_n148_ & new_nv452_;
  assign new_n_n41_ = ~new_n_n161_;
  assign new_n_n30_ = ~new_n_n150_;
  assign new_n_n19_ = ~new_n_n232_;
  assign new_n_n8_ = ~new_n_n221_;
  assign new_nv451_ = new_nv450_ & new_n_n271_;
  assign new_n_n40_ = ~new_n_n160_;
  assign new_n_n31_ = ~new_n_n151_;
  assign new_n_n18_ = ~new_n_n231_;
  assign new_n_n9_ = ~new_n_n222_;
  assign new_n_n39_ = ~new_n_n159_;
  assign new_n_n28_ = ~new_n_n241_;
  assign new_n_n21_ = ~new_n_n234_;
  assign new_n_n10_ = ~new_n_n223_;
  assign new_n_n38_ = ~new_n_n158_;
  assign new_n_n29_ = ~new_n_n242_;
  assign new_n_n20_ = ~new_n_n233_;
  assign new_n_n11_ = ~new_n_n224_;
  assign new_n_n67_ = ~new_n_n140_;
  assign new_n_n56_ = ~new_n_n176_;
  assign new_n_n45_ = ~new_n_n165_;
  assign new_n_n34_ = ~new_n_n154_;
  assign new_n_n23_ = ~new_n_n236_;
  assign new_n_n12_ = ~new_n_n225_;
  assign new_n_n66_ = ~new_n_n139_;
  assign new_n_n57_ = ~new_n_n177_;
  assign new_n_n44_ = ~new_n_n164_;
  assign new_n_n35_ = ~new_n_n155_;
  assign new_n_n22_ = ~new_n_n235_;
  assign new_n_n13_ = ~new_n_n226_;
  assign new_nv462_ = new_n_n140_ & new_nv453_ & new_n_n148_ & new_n_n272_;
  assign new_n_n68_ = new_nv460_ | new_nv480_ | new_nv467_ | new_nv482_;
  assign new_n_n43_ = ~new_n_n163_;
  assign new_n_n32_ = ~new_n_n152_;
  assign new_n_n25_ = ~new_n_n238_;
  assign new_n_n14_ = ~new_n_n227_;
  assign new_n_n73_ = new_nv455_ | new_nv475_ | new_nv462_ | new_nv482_;
  assign new_nv467_ = new_n_n135_ & new_nv453_ & new_n_n148_ & new_n_n272_;
  assign new_n_n42_ = ~new_n_n162_;
  assign new_n_n33_ = ~new_n_n153_;
  assign new_n_n24_ = ~new_n_n237_;
  assign new_n_n15_ = ~new_n_n228_;
  assign new_n_n74_ = new_nv474_ | new_nv461_ | new_nv454_;
  assign new_nv463_ = new_n_n139_ & new_nv453_ & new_n_n148_ & new_n_n272_;
  assign new_nv475_ = new_n_n67_ & new_n_n271_ & new_n_n148_ & new_n_n272_;
  assign new_n_n63_ = ~new_n_n136_;
  assign new_n_n52_ = ~new_n_n172_;
  assign new_n_n27_ = ~new_n_n240_;
  assign new_n_n16_ = ~new_n_n229_;
  assign new_nv461_ = new_n_n141_ & new_nv453_ & new_n_n148_ & new_n_n272_;
  assign new_n_n72_ = new_nv456_ | new_nv476_ | new_nv463_ | new_nv482_;
  assign new_nv474_ = new_n_n141_ & new_n_n271_ & new_n_n148_ & new_n_n272_;
  assign new_n_n62_ = ~new_n_n135_;
  assign new_n_n53_ = ~new_n_n173_;
  assign new_n_n26_ = ~new_n_n239_;
  assign new_n_n17_ = ~new_n_n230_;
  assign new_nv460_ = new_n_n142_ & new_nv453_ & new_n_n148_ & new_nv452_;
  assign new_nv464_ = new_n_n138_ & new_nv453_ & new_n_n148_ & new_n_n272_;
  assign new_nv477_ = new_n_n65_ & new_n_n271_ & new_n_n148_ & new_n_n272_;
  assign new_n_n65_ = ~new_n_n138_;
  assign new_n_n54_ = ~new_n_n174_;
  assign new_n_n47_ = ~new_n_n167_;
  assign new_n_n36_ = ~new_n_n156_;
  assign new_nv459_ = new_n_n143_ & new_nv453_ & new_n_n148_ & new_nv452_;
  assign new_n_n71_ = new_nv457_ | new_nv477_ | new_nv464_ | new_nv482_;
  assign new_nv476_ = new_n_n66_ & new_n_n271_ & new_n_n148_ & new_n_n272_;
  assign new_n_n64_ = ~new_n_n137_;
  assign new_n_n55_ = ~new_n_n175_;
  assign new_n_n46_ = ~new_n_n166_;
  assign new_n_n37_ = ~new_n_n157_;
endmodule


