// Benchmark "top" written by ABC on Fri Mar 31 12:08:23 2023

module top ( 
    pp, pa0, pq, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0, px,
    pi0, py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn,
    po,
    pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0  );
  input  pp, pa0, pq, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw,
    ph0, px, pi0, py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl,
    pm, pn, po;
  output pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0;
  wire new_np_, new_na0_, new_nq_, new_nr_, new_nc0_, new_ns_, new_nd0_,
    new_nt_, new_ne0_, new_nu_, new_nf0_, new_nv_, new_ng0_, new_nw_,
    new_nh0_, new_nx_, new_ni0_, new_ny_, new_nz_, new_na_, new_nb_,
    new_nc_, new_nd_, new_ne_, new_nf_, new_ng_, new_nh_, new_ni_, new_nj_,
    new_nk_, new_nl_, new_nm_, new_nn_, new_no_, new_np0_, new_nj1_,
    new_n_n435_, new_n_n426_, new_n_n418_, new_n_n411_, new_n_n402_,
    new_n_n395_, new_n_n386_, new_n_n376_, new_n_n367_, new_n_n360_,
    new_nc3_, new_n_n346_, new_n_n338_, new_n_n329_, new_n_n320_, new_nq3_,
    new_n_n300_, new_n_n293_, new_no4_, new_nt4_, new_n_n277_, new_n_n273_,
    new_nk5_, new_np5_, new_nh6_, new_n_n232_, new_n_n224_, new_nu6_,
    new_n_n210_, new_n_n201_, new_n_n193_, new_n_n158_, new_n_n147_,
    new_n_n136_, new_n_n125_, new_n_n114_, new_n_n103_, new_nk0_, new_no0_,
    new_n_n443_, new_nt1_, new_nx1_, new_n_n419_, new_n_n410_, new_nh2_,
    new_nn2_, new_n_n387_, new_n_n385_, new_n_n366_, new_n_n361_, new_nw5_,
    new_nf3_, new_n_n337_, new_n_n330_, new_n_n319_, new_n_n313_,
    new_n_n299_, new_n_n294_, new_np4_, new_ns4_, new_ny4_, new_nh5_,
    new_n_n264_, new_n_n258_, new_n_n245_, new_n_n231_, new_n_n225_,
    new_n_n218_, new_n_n211_, new_na7_, new_n_n194_, new_n_n157_,
    new_n_n148_, new_n_n135_, new_n_n126_, new_n_n113_, new_n_n104_,
    new_n_n442_, new_n_n433_, new_nw1_, new_n_n420_, new_n_n409_, new_ni2_,
    new_n_n396_, new_nq2_, new_nu2_, new_nz2_, new_n_n353_, new_ne3_,
    new_n_n336_, new_nl3_, new_nm3_, new_n_n314_, new_n_n298_, new_n_n292_,
    new_n_n291_, new_n_n284_, new_n_n276_, new_n_n271_, new_ni5_,
    new_n_n259_, new_n_n244_, new_n_n239_, new_nn6_, new_n_n217_,
    new_n_n208_, new_n_n203_, new_ne7_, new_nk7_, new_n_n167_, new_n_n134_,
    new_n_n123_, new_n_n116_, new_n_n105_, new_n_n441_, new_n_n434_,
    new_n_n427_, new_n_n421_, new_n_n408_, new_n_n401_, new_nm2_,
    new_n_n388_, new_nv2_, new_n_n359_, new_nb3_, new_n_n347_, new_n_n335_,
    new_n_n328_, new_n_n321_, new_np3_, new_n_n297_, new_nh4_, new_n_n290_,
    new_n_n285_, new_nz4_, new_n_n272_, new_nj5_, new_n_n260_, new_nd6_,
    new_ni6_, new_nk6_, new_n_n216_, new_n_n209_, new_n_n202_, new_n_n195_,
    new_n_n173_, new_nq7_, new_n_n133_, new_n_n124_, new_n_n115_,
    new_n_n106_, new_n_n450_, new_nr0_, new_n_n429_, new_nz1_, new_n_n382_,
    new_n_n374_, new_n_n348_, new_nj3_, new_n_n311_, new_nz3_, new_nb5_,
    new_n_n269_, new_n_n254_, new_nv5_, new_nv6_, new_ny6_, new_n_n198_,
    new_n_n190_, new_n_n181_, new_n_n132_, new_n_n121_, new_n_n110_,
    new_n_n99_, new_n_n9_, new_nl0_, new_n_n446_, new_n_n428_, new_ny1_,
    new_n_n381_, new_nt2_, new_n_n354_, new_n_n327_, new_nt3_, new_n_n304_,
    new_nc5_, new_n_n270_, new_nq5_, new_n_n249_, new_nw6_, new_n_n207_,
    new_n_n191_, new_ng7_, new_n_n182_, new_n_n131_, new_n_n122_,
    new_n_n109_, new_n_n100_, new_n_n452_, new_n_n447_, new_nh1_, new_ns1_,
    new_n_n384_, new_n_n375_, new_n_n362_, new_n_n318_, new_ns3_,
    new_n_n305_, new_n_n263_, new_n_n256_, new_n_n250_, new_n_n215_,
    new_n_n200_, new_n_n192_, new_n_n130_, new_n_n119_, new_n_n112_,
    new_n_n101_, new_n_n451_, new_nq0_, new_n_n444_, new_n_n436_,
    new_n_n383_, new_ns2_, new_n_n368_, new_nr3_, new_n_n312_, new_ny3_,
    new_nm5_, new_n_n257_, new_n_n255_, new_n_n206_, new_n_n199_, new_nf7_,
    new_n_n129_, new_n_n120_, new_n_n111_, new_n_n102_, new_nm0_,
    new_n_n445_, new_nk2_, new_n_n393_, new_n_n379_, new_n_n370_,
    new_n_n363_, new_n_n317_, new_n_n309_, new_n_n301_, new_nf4_, new_nn4_,
    new_ns5_, new_nx5_, new_ng6_, new_n_n234_, new_n_n226_, new_n_n187_,
    new_nj7_, new_no7_, new_n_n161_, new_n_n150_, new_n_n139_, new_n_n5_,
    new_nn0_, new_nf1_, new_n_n400_, new_n_n394_, new_n_n378_, new_n_n371_,
    new_n_n355_, new_n_n326_, new_n_n308_, new_na4_, new_ng4_, new_nm4_,
    new_nt5_, new_n_n246_, new_n_n241_, new_n_n235_, new_nt6_, new_ni7_,
    new_n_n178_, new_n_n169_, new_n_n162_, new_n_n149_, new_n_n140_,
    new_n_n6_, new_n_n449_, new_ne1_, new_n_n414_, new_n_n406_,
    new_n_n380_, new_n_n372_, new_n_n349_, new_n_n334_, new_nw3_,
    new_n_n302_, new_n_n287_, new_nw4_, new_nr5_, new_n_n247_, new_n_n240_,
    new_n_n228_, new_ns6_, new_n_n189_, new_n_n179_, new_n_n168_,
    new_n_n159_, new_n_n152_, new_n_n141_, new_n_n7_, new_n_n448_,
    new_ns0_, new_nd2_, new_n_n407_, new_nr2_, new_n_n373_, new_ni3_,
    new_n_n343_, new_n_n310_, new_n_n303_, new_n_n286_, new_nv4_,
    new_n_n253_, new_n_n248_, new_n_n233_, new_n_n227_, new_n_n222_,
    new_n_n188_, new_n_n180_, new_np7_, new_n_n160_, new_n_n151_,
    new_n_n142_, new_n_n8_, new_n_n440_, new_n_n431_, new_n_n423_,
    new_n_n415_, new_ne2_, new_n_n404_, new_n_n397_, new_n_n389_,
    new_n_n365_, new_n_n358_, new_n_n350_, new_n_n344_, new_n_n342_,
    new_n_n333_, new_n_n323_, new_no3_, new_n_n296_, new_nj4_, new_nr4_,
    new_n_n281_, new_nx4_, new_n_n274_, new_n_n266_, new_no5_, new_nu5_,
    new_ne6_, new_n_n237_, new_nm6_, new_n_n223_, new_n_n214_, new_n_n204_,
    new_n_n196_, new_n_n184_, new_n_n174_, new_n_n172_, new_n_n165_,
    new_n_n154_, new_n_n143_, new_n_n118_, new_n_n107_, new_n_n1_,
    new_n_n439_, new_n_n432_, new_n_n422_, new_n_n416_, new_n_n413_,
    new_n_n405_, new_nl2_, new_n_n390_, new_n_n364_, new_na3_, new_nd3_,
    new_nh3_, new_n_n341_, new_nk3_, new_n_n322_, new_nn3_, new_n_n295_,
    new_ni4_, new_n_n288_, new_n_n282_, new_n_n280_, new_n_n275_,
    new_n_n265_, new_nn5_, new_nc6_, new_n_n243_, new_n_n238_, new_n_n229_,
    new_nq6_, new_n_n221_, new_nz6_, new_n_n197_, new_n_n183_, new_n_n175_,
    new_nl7_, new_n_n166_, new_n_n153_, new_n_n144_, new_n_n117_,
    new_n_n108_, new_n_n2_, new_n_n438_, new_nu1_, new_n_n425_,
    new_n_n417_, new_n_n412_, new_ng2_, new_n_n399_, new_n_n391_,
    new_n_n377_, new_nw2_, new_n_n356_, new_n_n352_, new_ng3_, new_n_n340_,
    new_n_n331_, new_n_n325_, new_n_n315_, new_n_n307_, new_nc4_, new_nd4_,
    new_nl4_, new_n_n289_, new_n_n283_, new_n_n279_, new_ng5_, new_n_n268_,
    new_n_n261_, new_n_n252_, new_nb6_, new_n_n242_, new_n_n236_, new_nl6_,
    new_np6_, new_n_n220_, new_n_n212_, new_nb7_, new_n_n186_, new_n_n176_,
    new_n_n171_, new_n_n163_, new_n_n156_, new_n_n145_, new_n_n138_,
    new_n_n127_, new_n_n3_, new_n_n437_, new_n_n430_, new_n_n424_,
    new_na2_, new_nf2_, new_n_n403_, new_n_n398_, new_n_n392_, new_n_n369_,
    new_ny2_, new_n_n357_, new_n_n351_, new_n_n345_, new_n_n339_,
    new_n_n332_, new_n_n324_, new_n_n316_, new_n_n306_, new_nb4_, new_ne4_,
    new_nk4_, new_nq4_, new_nu4_, new_n_n278_, new_nf5_, new_n_n267_,
    new_n_n262_, new_n_n251_, new_ny5_, new_nf6_, new_nj6_, new_n_n230_,
    new_no6_, new_n_n219_, new_n_n213_, new_n_n205_, new_n_n185_,
    new_n_n177_, new_n_n170_, new_n_n164_, new_n_n155_, new_n_n146_,
    new_n_n137_, new_n_n128_, new_n_n4_, new_n_n93_, new_n_n82_,
    new_n_n71_, new_n_n61_, new_n_n50_, new_n_n94_, new_n_n81_, new_n_n72_,
    new_n_n60_, new_n_n51_, new_n_n95_, new_n_n80_, new_n_n69_, new_n_n63_,
    new_n_n52_, new_n_n96_, new_n_n79_, new_n_n70_, new_n_n62_, new_n_n53_,
    new_n_n0_, new_n_n97_, new_n_n43_, new_n_n32_, new_n_n21_, new_n_n10_,
    new_n_n98_, new_n_n42_, new_n_n33_, new_n_n20_, new_n_n11_, new_n_n41_,
    new_n_n30_, new_n_n23_, new_n_n12_, new_n_n40_, new_n_n31_, new_n_n22_,
    new_n_n13_, new_n_n68_, new_n_n58_, new_n_n47_, new_n_n36_, new_n_n25_,
    new_n_n14_, new_n_n67_, new_n_n59_, new_n_n46_, new_n_n37_, new_n_n24_,
    new_n_n15_, new_n_n88_, new_n_n77_, new_n_n45_, new_n_n34_, new_n_n27_,
    new_n_n16_, new_n_n87_, new_n_n78_, new_n_n44_, new_n_n35_, new_n_n26_,
    new_n_n17_, new_n_n89_, new_n_n86_, new_n_n75_, new_n_n64_, new_n_n54_,
    new_n_n29_, new_n_n18_, new_n_n90_, new_n_n85_, new_n_n76_, new_nj0_,
    new_n_n55_, new_n_n28_, new_n_n19_, new_n_n91_, new_n_n84_, new_n_n73_,
    new_n_n66_, new_n_n56_, new_n_n49_, new_n_n38_, new_n_n92_, new_n_n83_,
    new_n_n74_, new_n_n65_, new_n_n57_, new_n_n48_, new_n_n39_;
  assign new_np_ = pp;
  assign new_na0_ = pa0;
  assign new_nq_ = pq;
  assign new_nr_ = pr;
  assign new_nc0_ = pc0;
  assign new_ns_ = ps;
  assign new_nd0_ = pd0;
  assign new_nt_ = pt;
  assign new_ne0_ = pe0;
  assign new_nu_ = pu;
  assign new_nf0_ = pf0;
  assign new_nv_ = pv;
  assign new_ng0_ = pg0;
  assign new_nw_ = pw;
  assign new_nh0_ = ph0;
  assign new_nx_ = px;
  assign new_ni0_ = pi0;
  assign new_ny_ = py;
  assign pj0 = new_nj0_;
  assign new_nz_ = pz;
  assign pk0 = new_nk0_;
  assign pl0 = new_nl0_;
  assign pm0 = new_nm0_;
  assign pn0 = new_nn0_;
  assign po0 = new_no0_;
  assign pp0 = new_np0_;
  assign new_na_ = pa;
  assign pq0 = new_nq0_;
  assign new_nb_ = pb;
  assign pr0 = new_nr0_;
  assign new_nc_ = pc;
  assign ps0 = new_ns0_;
  assign new_nd_ = pd;
  assign new_ne_ = pe;
  assign new_nf_ = pf;
  assign new_ng_ = pg;
  assign new_nh_ = ph;
  assign new_ni_ = pi;
  assign new_nj_ = pj;
  assign new_nk_ = pk;
  assign new_nl_ = pl;
  assign new_nm_ = pm;
  assign new_nn_ = pn;
  assign new_no_ = po;
  assign new_np0_ = new_nb_ & new_n_n8_ & new_n_n7_;
  assign new_nj1_ = new_n_n438_ | new_n_n437_ | new_n_n443_ | new_n_n436_ | new_n_n442_ | new_n_n441_ | new_n_n440_ | new_n_n439_;
  assign new_n_n435_ = new_n_n129_ & new_n_n133_;
  assign new_n_n426_ = new_n_n18_ & new_n_n161_;
  assign new_n_n418_ = new_nt_ & new_nq_ & new_n_n20_;
  assign new_n_n411_ = new_n_n133_ & new_n_n131_ & new_n_n23_;
  assign new_n_n402_ = new_n_n25_ & new_n_n133_;
  assign new_n_n395_ = new_n_n107_ & new_n_n49_;
  assign new_n_n386_ = new_nu_ & new_nq_ & new_ns_;
  assign new_n_n376_ = new_nr_ & new_nt_ & new_n_n32_;
  assign new_n_n367_ = new_n_n33_ & new_n_n35_ & new_n_n34_;
  assign new_n_n360_ = new_np_ & new_nv_ & new_n_n40_;
  assign new_nc3_ = new_n_n351_ | new_nw5_ | new_n_n350_ | new_n_n352_;
  assign new_n_n346_ = new_n_n44_ & new_nr_;
  assign new_n_n338_ = new_n_n131_ & new_n_n63_;
  assign new_n_n329_ = new_n_n140_ & new_n_n52_ & new_n_n47_;
  assign new_n_n320_ = new_nt_ & new_nx_ & new_nr_;
  assign new_nq3_ = new_n_n121_ & new_nf0_ & new_n_n59_;
  assign new_n_n300_ = new_n_n122_ & new_nq_ & new_n_n74_;
  assign new_n_n293_ = new_nr_ & new_nt_ & new_n_n76_;
  assign new_no4_ = new_n_n124_ | new_np_ | new_n_n119_;
  assign new_nt4_ = new_nt_ & new_ns_ & new_n_n140_;
  assign new_n_n277_ = new_nf0_ & new_n_n91_ & new_n_n90_;
  assign new_n_n273_ = new_n_n94_ & new_ni0_ & new_n_n96_;
  assign new_nk5_ = new_n_n263_ | new_n_n264_;
  assign new_np5_ = new_n_n255_ | new_n_n257_ | new_n_n254_ | new_n_n256_;
  assign new_nh6_ = new_nq_ | new_n_n142_ | new_n_n130_;
  assign new_n_n232_ = new_n_n140_ & new_n_n134_;
  assign new_n_n224_ = new_n_n143_ & new_n_n140_;
  assign new_nu6_ = new_n_n218_ | new_n_n217_ | new_n_n216_;
  assign new_n_n210_ = new_n_n149_ & new_nd_ & new_n_n147_;
  assign new_n_n201_ = new_n_n152_ & new_nd_;
  assign new_n_n193_ = new_ne_ & new_nd_;
  assign new_n_n158_ = ~new_no7_;
  assign new_n_n147_ = ~new_nk7_;
  assign new_n_n136_ = ~new_nm4_;
  assign new_n_n125_ = ~new_nl6_;
  assign new_n_n114_ = ~new_nt5_;
  assign new_n_n103_ = ~new_nb6_;
  assign new_nk0_ = new_n_n452_ | new_n_n451_ | new_n_n450_;
  assign new_no0_ = new_nb_ & new_n_n8_ & new_n_n6_;
  assign new_n_n443_ = new_np_ & new_nq_ & new_nr_;
  assign new_nt1_ = new_n_n435_ | new_n_n434_ | new_n_n433_ | new_n_n432_ | new_n_n430_ | new_n_n400_ | new_n_n431_;
  assign new_nx1_ = new_n_n423_ | new_n_n425_ | new_n_n422_ | new_n_n424_;
  assign new_n_n419_ = new_ny_ & new_nq_ & new_n_n20_;
  assign new_n_n410_ = new_n_n22_ & new_n_n131_ & new_n_n23_;
  assign new_nh2_ = new_n_n401_ | new_n_n402_;
  assign new_nn2_ = new_n_n390_ | new_n_n389_ | new_nj5_ | new_n_n388_ | new_n_n394_ | new_n_n393_ | new_n_n392_ | new_n_n391_;
  assign new_n_n387_ = new_np_ & new_nq_ & new_ns_;
  assign new_n_n385_ = new_np_ & new_nv_ & new_ns_;
  assign new_n_n366_ = new_n_n36_ & new_n_n35_ & new_n_n34_;
  assign new_n_n361_ = new_nu_ & new_nq_ & new_n_n40_;
  assign new_nw5_ = new_ns_ & new_nt_;
  assign new_nf3_ = new_n_n43_ | new_n_n346_ | new_n_n345_;
  assign new_n_n337_ = new_n_n143_ & new_n_n46_ & new_n_n133_;
  assign new_n_n330_ = new_n_n62_ & new_n_n52_ & new_n_n47_;
  assign new_n_n319_ = new_ny_ & new_nx_ & new_nr_;
  assign new_n_n313_ = new_n_n162_ & new_n_n58_ & new_n_n57_;
  assign new_n_n299_ = new_n_n131_ & new_nq_ & new_n_n74_;
  assign new_n_n294_ = new_n_n76_ & new_ns_;
  assign new_np4_ = new_n_n289_ | new_n_n82_;
  assign new_ns4_ = new_nq_ & new_np_ & new_nm_;
  assign new_ny4_ = new_nt_ | new_n_n92_ | new_n_n276_;
  assign new_nh5_ = new_n_n268_ | new_n_n267_ | new_n_n266_ | new_n_n265_ | new_n_n272_ | new_n_n270_ | new_n_n269_ | new_n_n271_ | new_n_n273_;
  assign new_n_n264_ = new_ne0_ & new_n_n103_ & new_n_n115_;
  assign new_n_n258_ = new_n_n110_ & new_n_n109_ & new_n_n108_;
  assign new_n_n245_ = new_n_n130_ & new_n_n124_;
  assign new_n_n231_ = new_n_n134_ & new_ns_ & new_nt_;
  assign new_n_n225_ = new_n_n139_ & new_n_n140_;
  assign new_n_n218_ = new_n_n145_ & new_n_n161_;
  assign new_n_n211_ = new_nc_ & new_nd_ & new_n_n147_;
  assign new_na7_ = new_n_n200_ | new_n_n199_ | new_n_n198_;
  assign new_n_n194_ = new_nh_ & new_nd_;
  assign new_n_n157_ = ~new_np7_;
  assign new_n_n148_ = ~new_nj7_;
  assign new_n_n135_ = ~new_nn4_;
  assign new_n_n126_ = ~new_nj6_;
  assign new_n_n113_ = ~new_nx5_;
  assign new_n_n104_ = ~new_ne6_;
  assign new_n_n442_ = new_nu_ & new_nq_ & new_nr_;
  assign new_n_n433_ = new_n_n16_ & new_nd0_;
  assign new_nw1_ = new_n_n426_ | new_n_n427_;
  assign new_n_n420_ = new_nt_ & new_nv_ & new_n_n20_;
  assign new_n_n409_ = new_n_n36_ & new_n_n131_ & new_n_n23_;
  assign new_ni2_ = new_ne0_ & new_n_n161_ & new_n_n27_;
  assign new_n_n396_ = new_n_n140_ & new_n_n61_;
  assign new_nq2_ = new_n_n382_ | new_n_n381_ | new_n_n387_ | new_n_n380_ | new_n_n386_ | new_n_n385_ | new_n_n384_ | new_n_n383_;
  assign new_nu2_ = new_n_n122_ & new_ne0_ & new_nd0_;
  assign new_nz2_ = new_n_n131_ | new_n_n129_ | new_n_n133_;
  assign new_n_n353_ = new_n_n42_ & new_n_n48_ & new_n_n41_;
  assign new_ne3_ = new_ne0_ & new_nd0_ & new_nc0_;
  assign new_n_n336_ = new_n_n143_ & new_n_n46_ & new_n_n129_;
  assign new_nl3_ = new_n_n326_ | new_n_n324_ | new_n_n323_ | new_n_n322_ | new_n_n325_ | new_n_n327_;
  assign new_nm3_ = new_n_n317_ | new_n_n316_ | new_ns5_ | new_n_n315_ | new_n_n321_ | new_n_n320_ | new_n_n319_ | new_n_n318_;
  assign new_n_n314_ = new_n_n161_ & new_n_n58_ & new_n_n57_;
  assign new_n_n298_ = new_n_n91_ & new_nq_ & new_n_n74_;
  assign new_n_n292_ = new_n_n140_ & new_n_n143_;
  assign new_n_n291_ = new_nt_ & new_n_n80_;
  assign new_n_n284_ = new_n_n88_ & new_n_n87_ & new_n_n86_;
  assign new_n_n276_ = new_n_n122_ & new_n_n129_ & new_n_n133_;
  assign new_n_n271_ = new_n_n98_ & new_ni0_ & new_n_n96_;
  assign new_ni5_ = new_n_n107_ & new_nk_ & new_n_n99_;
  assign new_n_n259_ = new_n_n107_ & new_n_n109_ & new_n_n108_;
  assign new_n_n244_ = new_n_n125_ & new_nq_;
  assign new_n_n239_ = new_n_n143_ & new_n_n139_;
  assign new_nn6_ = new_n_n138_ | new_n_n225_ | new_n_n224_;
  assign new_n_n217_ = new_nc_ & new_n_n161_;
  assign new_n_n208_ = new_nc_ & new_n_n148_ & new_n_n147_;
  assign new_n_n203_ = new_n_n152_ & new_n_n164_;
  assign new_ne7_ = new_n_n194_ | new_n_n193_ | new_n_n187_;
  assign new_nk7_ = new_n_n172_ | new_n_n173_;
  assign new_n_n167_ = new_nd_ & new_n_n164_ & new_ne_;
  assign new_n_n134_ = ~new_nm_;
  assign new_n_n123_ = ~new_nm6_;
  assign new_n_n116_ = ~new_nu5_;
  assign new_n_n105_ = ~new_nd6_;
  assign new_n_n441_ = new_np_ & new_nv_ & new_nr_;
  assign new_n_n434_ = new_n_n16_ & new_n_n133_;
  assign new_n_n427_ = new_n_n18_ & new_n_n162_;
  assign new_n_n421_ = new_ny_ & new_nv_ & new_n_n20_;
  assign new_n_n408_ = new_n_n133_ & new_nc_ & new_n_n23_;
  assign new_n_n401_ = new_n_n26_ & new_n_n129_;
  assign new_nm2_ = new_n_n31_ | new_ng3_ | new_n_n395_;
  assign new_n_n388_ = new_nx_ & new_nw_ & new_nv_;
  assign new_nv2_ = new_n_n37_ | new_n_n365_ | new_n_n364_;
  assign new_n_n359_ = new_nu_ & new_nv_ & new_n_n40_;
  assign new_nb3_ = new_nt_ | new_ny_;
  assign new_n_n347_ = new_nw_ & new_nt_ & new_nx_;
  assign new_n_n335_ = new_n_n143_ & new_n_n46_ & new_n_n131_;
  assign new_n_n328_ = new_n_n48_ & new_n_n52_ & new_n_n47_;
  assign new_n_n321_ = new_ny_ & new_ns_ & new_nr_;
  assign new_np3_ = new_n_n313_ | new_n_n314_;
  assign new_n_n297_ = new_n_n122_ & new_n_n118_ & new_n_n74_;
  assign new_nh4_ = new_n_n121_ | new_n_n77_ | new_n_n292_;
  assign new_n_n290_ = new_ns_ & new_n_n81_;
  assign new_n_n285_ = new_n_n85_ & new_n_n87_ & new_n_n86_;
  assign new_nz4_ = new_np_ & new_no_ & new_n_n93_;
  assign new_n_n272_ = new_n_n95_ & new_ni0_ & new_n_n96_;
  assign new_nj5_ = new_ns_ & new_nr_ & new_nq_;
  assign new_n_n260_ = new_np_ & new_n_n110_ & new_n_n108_;
  assign new_nd6_ = new_nf0_ | new_ng0_;
  assign new_ni6_ = new_n_n239_ | new_n_n238_ | new_n_n237_;
  assign new_nk6_ = new_n_n224_ | new_n_n232_ | new_n_n231_ | new_n_n225_;
  assign new_n_n216_ = new_nc_ & new_n_n145_;
  assign new_n_n209_ = new_n_n159_ & new_n_n148_ & new_n_n147_;
  assign new_n_n202_ = new_n_n152_ & new_n_n163_;
  assign new_n_n195_ = new_n_n154_ & new_nd_;
  assign new_n_n173_ = new_n_n160_ & new_n_n164_;
  assign new_nq7_ = new_n_n166_ | new_n_n167_;
  assign new_n_n133_ = ~new_nc0_;
  assign new_n_n124_ = ~new_nq_;
  assign new_n_n115_ = ~new_nf5_;
  assign new_n_n106_ = ~new_no5_;
  assign new_n_n450_ = new_n_n0_ & new_n_n162_;
  assign new_nr0_ = new_n_n58_ & new_na_ & new_n_n12_;
  assign new_n_n429_ = new_n_n26_ & new_n_n162_;
  assign new_nz1_ = new_n_n419_ | new_n_n421_ | new_n_n418_ | new_n_n420_;
  assign new_n_n382_ = new_nu_ & new_nq_ & new_nx_;
  assign new_n_n374_ = new_n_n133_ & new_n_n122_ & new_n_n34_;
  assign new_n_n348_ = new_nw_ & new_ny_ & new_nx_;
  assign new_nj3_ = new_n_n344_ | new_n_n334_ | new_n_n412_;
  assign new_n_n311_ = new_n_n60_ & new_nt_;
  assign new_nz3_ = new_n_n70_ | new_n_n303_ | new_n_n302_;
  assign new_nb5_ = new_n_n139_ | new_n_n140_ | new_n_n124_;
  assign new_n_n269_ = new_n_n95_ & new_n_n107_ & new_n_n96_;
  assign new_n_n254_ = new_n_n113_ & new_n_n112_ & new_n_n111_;
  assign new_nv5_ = new_n_n248_ | new_n_n247_ | new_n_n246_;
  assign new_nv6_ = new_n_n146_ | new_nj_;
  assign new_ny6_ = new_n_n206_ | new_n_n205_ | new_n_n204_;
  assign new_n_n198_ = new_n_n153_ & new_n_n161_;
  assign new_n_n190_ = new_n_n155_ & new_n_n161_;
  assign new_n_n181_ = new_n_n158_ & new_ne_ & new_n_n156_;
  assign new_n_n132_ = ~new_nk6_;
  assign new_n_n121_ = ~new_ng0_;
  assign new_n_n110_ = ~new_np5_;
  assign new_n_n99_ = ~new_ns6_;
  assign new_n_n9_ = ~new_nl3_;
  assign new_nl0_ = new_n_n448_ | new_n_n449_;
  assign new_n_n446_ = new_nu_ & new_nq_ & new_n_n11_;
  assign new_n_n428_ = new_n_n17_ & new_n_n161_;
  assign new_ny1_ = new_n_n413_ | new_n_n344_ | new_n_n334_;
  assign new_n_n381_ = new_np_ & new_nv_ & new_nx_;
  assign new_nt2_ = new_n_n369_ | new_n_n368_ | new_n_n367_ | new_n_n366_ | new_n_n373_ | new_n_n371_ | new_n_n370_ | new_n_n372_ | new_n_n374_;
  assign new_n_n354_ = new_n_n139_ & new_n_n48_ & new_n_n41_;
  assign new_n_n327_ = new_n_n62_ & new_n_n121_ & new_n_n50_;
  assign new_nt3_ = new_n_n61_ | new_n_n62_ | new_n_n334_;
  assign new_n_n304_ = new_n_n118_ & new_n_n69_ & new_n_n68_;
  assign new_nc5_ = new_n_n274_ | new_n_n275_;
  assign new_n_n270_ = new_n_n94_ & new_n_n107_ & new_n_n96_;
  assign new_nq5_ = new_n_n140_ | new_n_n124_ | new_n_n120_;
  assign new_n_n249_ = new_nq_ & new_n_n119_ & new_n_n118_;
  assign new_nw6_ = new_n_n210_ | new_n_n209_ | new_n_n208_ | new_n_n207_ | new_n_n214_ | new_n_n212_ | new_n_n211_ | new_n_n213_ | new_n_n215_;
  assign new_n_n207_ = new_n_n149_ & new_n_n148_ & new_n_n147_;
  assign new_n_n191_ = new_n_n155_ & new_ne_;
  assign new_ng7_ = new_n_n189_ | new_n_n188_ | new_n_n187_;
  assign new_n_n182_ = new_nd_ & new_ne_ & new_n_n156_;
  assign new_n_n131_ = ~new_ne0_;
  assign new_n_n122_ = ~new_nf0_;
  assign new_n_n109_ = ~new_nq5_;
  assign new_n_n100_ = ~new_nq6_;
  assign new_n_n452_ = new_n_n0_ & new_nj0_;
  assign new_n_n447_ = new_n_n10_ & new_np_;
  assign new_nh1_ = new_n_n15_ | new_n_n444_ | new_ng3_;
  assign new_ns1_ = new_n_n55_ | new_na0_;
  assign new_n_n384_ = new_nu_ & new_nv_ & new_ns_;
  assign new_n_n375_ = new_n_n62_ & new_n_n124_;
  assign new_n_n362_ = new_np_ & new_nq_ & new_n_n40_;
  assign new_n_n318_ = new_nt_ & new_ns_ & new_nw_;
  assign new_ns3_ = new_n_n311_ | new_n_n312_;
  assign new_n_n305_ = new_n_n118_ & new_n_n67_ & new_n_n69_;
  assign new_n_n263_ = new_n_n121_ & new_n_n122_ & new_n_n100_;
  assign new_n_n256_ = new_n_n113_ & new_nr_ & new_n_n111_;
  assign new_n_n250_ = new_n_n140_ & new_n_n139_;
  assign new_n_n215_ = new_n_n159_ & new_n_n165_ & new_n_n147_;
  assign new_n_n200_ = new_n_n153_ & new_n_n164_;
  assign new_n_n192_ = new_n_n155_ & new_nh_;
  assign new_n_n130_ = ~new_ns5_;
  assign new_n_n119_ = ~new_nk_;
  assign new_n_n112_ = ~new_ny5_;
  assign new_n_n101_ = ~new_nf6_;
  assign new_n_n451_ = new_n_n0_ & new_nd_;
  assign new_nq0_ = new_n_n9_ | new_n_n447_ | new_n_n446_;
  assign new_n_n444_ = new_n_n139_ & new_n_n63_;
  assign new_n_n436_ = new_nu_ & new_nv_ & new_nw_;
  assign new_n_n383_ = new_np_ & new_nq_ & new_nx_;
  assign new_ns2_ = new_n_n413_ | new_n_n375_ | new_n_n334_;
  assign new_n_n368_ = new_n_n133_ & new_n_n35_ & new_n_n34_;
  assign new_nr3_ = new_ne0_ & new_nf0_;
  assign new_n_n312_ = new_n_n60_ & new_ny_;
  assign new_ny3_ = new_n_n66_ | new_n_n305_ | new_n_n304_;
  assign new_nm5_ = new_n_n101_ | new_n_n262_ | new_n_n261_;
  assign new_n_n257_ = new_nq_ & new_nr_ & new_n_n111_;
  assign new_n_n255_ = new_nq_ & new_n_n112_ & new_n_n111_;
  assign new_n_n206_ = new_n_n151_ & new_n_n162_;
  assign new_n_n199_ = new_n_n153_ & new_n_n163_;
  assign new_nf7_ = new_n_n192_ | new_n_n191_ | new_n_n190_;
  assign new_n_n129_ = ~new_nd0_;
  assign new_n_n120_ = ~new_nw5_;
  assign new_n_n111_ = ~new_ni6_;
  assign new_n_n102_ = ~new_nc6_;
  assign new_nm0_ = new_nb_ & new_n_n4_ & new_n_n3_;
  assign new_n_n445_ = new_nd_ & new_nc_;
  assign new_nk2_ = new_n_n398_ | new_n_n400_ | new_n_n397_ | new_n_n399_;
  assign new_n_n393_ = new_ns_ & new_nw_ & new_nq_;
  assign new_n_n379_ = new_nw_ & new_ny_ & new_n_n32_;
  assign new_n_n370_ = new_n_n33_ & new_nc_ & new_n_n34_;
  assign new_n_n363_ = new_n_n40_ & new_n_n59_;
  assign new_n_n317_ = new_ny_ & new_ns_ & new_nw_;
  assign new_n_n309_ = new_n_n65_ & new_nj0_;
  assign new_n_n301_ = new_n_n73_ & new_n_n124_;
  assign new_nf4_ = new_n_n75_ | new_n_n275_ | new_n_n274_;
  assign new_nn4_ = new_n_n291_ | new_n_n290_ | new_nw5_;
  assign new_ns5_ = new_nt_ & new_ns_ & new_nr_;
  assign new_nx5_ = new_n_n140_ | new_nl_ | new_n_n120_;
  assign new_ng6_ = new_n_n240_ | new_n_n241_;
  assign new_n_n234_ = new_n_n131_ & new_ns_ & new_n_n132_;
  assign new_n_n226_ = new_nc0_ & new_ns_ & new_n_n137_;
  assign new_n_n187_ = new_ne_ & new_nh_;
  assign new_nj7_ = new_n_n175_ | new_n_n177_ | new_n_n174_ | new_n_n176_;
  assign new_no7_ = new_n_n168_ | new_n_n169_;
  assign new_n_n161_ = ~new_nd_;
  assign new_n_n150_ = ~new_na7_;
  assign new_n_n139_ = ~new_ns_;
  assign new_n_n5_ = ~new_nt1_;
  assign new_nn0_ = new_nb_ & new_n_n8_ & new_n_n5_;
  assign new_nf1_ = new_n_n445_ | new_n_n14_;
  assign new_n_n400_ = new_nd0_ & new_nc0_;
  assign new_n_n394_ = new_nx_ & new_nr_ & new_nq_;
  assign new_n_n378_ = new_nr_ & new_ny_ & new_n_n32_;
  assign new_n_n371_ = new_n_n133_ & new_nc_ & new_n_n34_;
  assign new_n_n355_ = new_n_n61_ & new_n_n48_ & new_n_n41_;
  assign new_n_n326_ = new_n_n49_ & new_n_n121_ & new_n_n50_;
  assign new_n_n308_ = new_n_n64_ & new_n_n121_;
  assign new_na4_ = new_n_n135_ | new_n_n301_ | new_n_n230_;
  assign new_ng4_ = new_n_n293_ | new_n_n294_;
  assign new_nm4_ = new_nt_ & new_ns_ & new_n_n134_;
  assign new_nt5_ = new_n_n251_ | new_n_n252_;
  assign new_n_n246_ = new_nd0_ & new_ne0_ & new_nf0_;
  assign new_n_n241_ = new_n_n128_ & new_n_n131_;
  assign new_n_n235_ = new_n_n133_ & new_nt_ & new_n_n132_;
  assign new_nt6_ = new_n_n221_ | new_n_n220_ | new_n_n219_;
  assign new_ni7_ = new_n_n181_ | new_n_n180_ | new_n_n179_ | new_n_n178_ | new_n_n185_ | new_n_n183_ | new_n_n182_ | new_n_n184_ | new_n_n186_;
  assign new_n_n178_ = new_n_n158_ & new_n_n157_ & new_n_n156_;
  assign new_n_n169_ = new_nh_ & new_ne_;
  assign new_n_n162_ = ~new_nc_;
  assign new_n_n149_ = ~new_ni7_;
  assign new_n_n140_ = ~new_nr_;
  assign new_n_n6_ = ~new_nf2_;
  assign new_n_n449_ = new_n_n54_ & new_n_n2_ & new_n_n1_;
  assign new_ne1_ = new_nc0_ | new_na0_ | new_n_n55_;
  assign new_n_n414_ = new_nt_ & new_np_ & new_n_n21_;
  assign new_n_n406_ = new_n_n36_ & new_nc_ & new_n_n23_;
  assign new_n_n380_ = new_nu_ & new_nv_ & new_nx_;
  assign new_n_n372_ = new_n_n36_ & new_n_n122_ & new_n_n34_;
  assign new_n_n349_ = new_nc0_ & new_nd0_ & new_ne0_;
  assign new_n_n334_ = new_n_n63_ & new_n_n139_;
  assign new_nw3_ = new_n_n309_ | new_n_n307_ | new_n_n306_ | new_n_n308_ | new_n_n310_;
  assign new_n_n302_ = new_n_n72_ & new_n_n107_;
  assign new_n_n287_ = new_n_n85_ & new_n_n84_ & new_n_n86_;
  assign new_nw4_ = new_nt_ & new_n_n139_ & new_nr_;
  assign new_nr5_ = new_n_n114_ | new_n_n245_ | new_n_n253_;
  assign new_n_n247_ = new_nc0_ & new_ne0_ & new_nf0_;
  assign new_n_n240_ = new_n_n133_ & new_n_n129_ & new_n_n128_;
  assign new_n_n228_ = new_nc0_ & new_nt_ & new_n_n137_;
  assign new_ns6_ = new_n_n143_ | new_ni0_;
  assign new_n_n189_ = new_nh_ & new_n_n161_;
  assign new_n_n179_ = new_nd_ & new_n_n157_ & new_n_n156_;
  assign new_n_n168_ = new_n_n164_ & new_n_n163_;
  assign new_n_n159_ = ~new_ng_;
  assign new_n_n152_ = ~new_nf7_;
  assign new_n_n141_ = ~new_np6_;
  assign new_n_n7_ = ~new_nt2_;
  assign new_n_n448_ = new_nb_ & new_n_n2_ & new_ny6_;
  assign new_ns0_ = new_n_n58_ & new_na_ & new_n_n13_;
  assign new_nd2_ = new_n_n334_ | new_n_n375_ | new_n_n412_;
  assign new_n_n407_ = new_n_n22_ & new_nc_ & new_n_n23_;
  assign new_nr2_ = new_n_n377_ | new_n_n379_ | new_n_n376_ | new_n_n378_;
  assign new_n_n373_ = new_n_n33_ & new_n_n122_ & new_n_n34_;
  assign new_ni3_ = new_n_n338_ | new_n_n337_ | new_n_n336_ | new_n_n335_ | new_n_n342_ | new_n_n340_ | new_n_n339_ | new_n_n341_ | new_n_n343_;
  assign new_n_n343_ = new_n_n133_ & new_n_n61_;
  assign new_n_n310_ = new_nj0_ & new_n_n121_;
  assign new_n_n303_ = new_n_n71_ & new_np_;
  assign new_n_n286_ = new_n_n88_ & new_n_n84_ & new_n_n86_;
  assign new_nv4_ = new_nq_ & new_np_ & new_nn_;
  assign new_n_n253_ = new_n_n121_ & new_ne0_ & new_n_n115_;
  assign new_n_n248_ = new_n_n121_ & new_n_n122_;
  assign new_n_n233_ = new_n_n133_ & new_ns_ & new_n_n132_;
  assign new_n_n227_ = new_nd0_ & new_ns_ & new_n_n137_;
  assign new_n_n222_ = new_ne0_ & new_nd0_;
  assign new_n_n188_ = new_ne_ & new_n_n161_;
  assign new_n_n180_ = new_n_n165_ & new_n_n157_ & new_n_n156_;
  assign new_np7_ = new_nd_ | new_n_n165_;
  assign new_n_n160_ = ~new_nl7_;
  assign new_n_n151_ = ~new_nz6_;
  assign new_n_n142_ = ~new_nl_;
  assign new_n_n8_ = ~new_ns1_;
  assign new_n_n440_ = new_nu_ & new_nv_ & new_nr_;
  assign new_n_n431_ = new_n_n36_ & new_n_n129_;
  assign new_n_n423_ = new_nw_ & new_nq_ & new_n_n19_;
  assign new_n_n415_ = new_ny_ & new_np_ & new_n_n21_;
  assign new_ne2_ = new_n_n413_ | new_n_n334_ | new_n_n412_;
  assign new_n_n404_ = new_n_n22_ & new_n_n24_ & new_n_n23_;
  assign new_n_n397_ = new_n_n28_ & new_n_n29_;
  assign new_n_n389_ = new_ns_ & new_nw_ & new_nv_;
  assign new_n_n365_ = new_n_n107_ & new_n_n49_ & new_n_n38_;
  assign new_n_n358_ = new_n_n61_ & new_n_n140_ & new_n_n41_;
  assign new_n_n350_ = new_nx_ & new_ny_;
  assign new_n_n344_ = new_n_n46_ & new_n_n143_;
  assign new_n_n342_ = new_n_n133_ & new_n_n63_;
  assign new_n_n333_ = new_n_n62_ & new_n_n124_ & new_n_n47_;
  assign new_n_n323_ = new_n_n49_ & new_n_n51_ & new_n_n50_;
  assign new_no3_ = new_n_n54_ | new_n_n55_ | new_n_n56_;
  assign new_n_n296_ = new_n_n131_ & new_n_n118_ & new_n_n74_;
  assign new_nj4_ = new_nr_ & new_nq_ & new_n_n119_;
  assign new_nr4_ = new_n_n287_ | new_n_n285_ | new_n_n284_ | new_n_n286_ | new_n_n288_;
  assign new_n_n281_ = new_n_n89_ & new_n_n91_;
  assign new_nx4_ = new_n_n278_ | new_n_n280_ | new_n_n277_ | new_n_n279_;
  assign new_n_n274_ = new_n_n133_ & new_n_n129_ & new_n_n122_;
  assign new_n_n266_ = new_n_n95_ & new_n_n97_ & new_n_n96_;
  assign new_no5_ = new_n_n260_ | new_n_n259_ | new_n_n258_;
  assign new_nu5_ = new_n_n117_ | new_n_n250_ | new_n_n249_;
  assign new_ne6_ = new_n_n126_ | new_n_n243_ | new_n_n242_;
  assign new_n_n237_ = new_nn_ & new_n_n139_;
  assign new_nm6_ = new_n_n227_ | new_n_n229_ | new_n_n226_ | new_n_n228_;
  assign new_n_n223_ = new_ne0_ & new_nc0_;
  assign new_n_n214_ = new_nc_ & new_n_n165_ & new_n_n147_;
  assign new_n_n204_ = new_n_n150_ & new_n_n151_;
  assign new_n_n196_ = new_n_n154_ & new_ne_;
  assign new_n_n184_ = new_n_n158_ & new_n_n164_ & new_n_n156_;
  assign new_n_n174_ = new_n_n163_ & new_n_n159_ & new_n_n164_;
  assign new_n_n172_ = new_n_n160_ & new_n_n163_;
  assign new_n_n165_ = ~new_nf_;
  assign new_n_n154_ = ~new_ne7_;
  assign new_n_n143_ = ~new_nt_;
  assign new_n_n118_ = ~new_ne4_;
  assign new_n_n107_ = ~new_np_;
  assign new_n_n1_ = ~new_nw6_;
  assign new_n_n439_ = new_np_ & new_nq_ & new_nw_;
  assign new_n_n432_ = new_n_n36_ & new_nc0_;
  assign new_n_n422_ = new_nr_ & new_nq_ & new_n_n19_;
  assign new_n_n416_ = new_nt_ & new_nu_ & new_n_n21_;
  assign new_n_n413_ = new_n_n49_ & new_n_n107_;
  assign new_n_n405_ = new_n_n133_ & new_n_n24_ & new_n_n23_;
  assign new_nl2_ = new_n_n30_ | new_n_n396_ | new_ng3_;
  assign new_n_n390_ = new_nx_ & new_nr_ & new_nv_;
  assign new_n_n364_ = new_n_n124_ & new_n_n62_ & new_n_n38_;
  assign new_na3_ = new_n_n357_ | new_n_n355_ | new_n_n354_ | new_n_n353_ | new_n_n356_ | new_n_n358_;
  assign new_nd3_ = new_n_n349_ | new_n_n348_ | new_n_n347_;
  assign new_nh3_ = new_n_n334_ | new_n_n344_;
  assign new_n_n341_ = new_n_n129_ & new_n_n61_;
  assign new_nk3_ = new_n_n332_ | new_n_n330_ | new_n_n329_ | new_n_n328_ | new_n_n331_ | new_n_n333_;
  assign new_n_n322_ = new_n_n52_ & new_n_n51_ & new_n_n50_;
  assign new_nn3_ = new_n_n129_ | new_n_n133_ | new_n_n53_;
  assign new_n_n295_ = new_n_n91_ & new_n_n118_ & new_n_n74_;
  assign new_ni4_ = new_n_n143_ | new_n_n139_ | new_n_n78_;
  assign new_n_n288_ = new_n_n86_ & new_n_n83_;
  assign new_n_n282_ = new_n_n89_ & new_n_n131_;
  assign new_n_n280_ = new_n_n131_ & new_nf0_ & new_n_n90_;
  assign new_n_n275_ = new_n_n122_ & new_n_n131_;
  assign new_n_n265_ = new_n_n98_ & new_n_n97_ & new_n_n96_;
  assign new_nn5_ = new_n_n106_ & new_ni0_;
  assign new_nc6_ = new_n_n123_ | new_n_n245_ | new_n_n244_;
  assign new_n_n243_ = new_n_n111_ & new_nr_;
  assign new_n_n238_ = new_no_ & new_n_n143_;
  assign new_n_n229_ = new_nd0_ & new_nt_ & new_n_n137_;
  assign new_nq6_ = new_n_n222_ | new_n_n223_;
  assign new_n_n221_ = new_n_n144_ & new_nh0_;
  assign new_nz6_ = new_n_n203_ | new_n_n202_ | new_n_n201_;
  assign new_n_n197_ = new_n_n154_ & new_nh_;
  assign new_n_n183_ = new_n_n165_ & new_ne_ & new_n_n156_;
  assign new_n_n175_ = new_nc_ & new_n_n163_ & new_n_n164_;
  assign new_nl7_ = new_n_n171_ | new_n_n168_ | new_n_n170_;
  assign new_n_n166_ = new_n_n165_ & new_n_n164_ & new_ne_;
  assign new_n_n153_ = ~new_nb7_;
  assign new_n_n144_ = ~new_nu6_;
  assign new_n_n117_ = ~new_nv5_;
  assign new_n_n108_ = ~new_nr5_;
  assign new_n_n2_ = ~new_nv6_;
  assign new_n_n438_ = new_nu_ & new_nq_ & new_nw_;
  assign new_nu1_ = new_n_n428_ | new_n_n429_;
  assign new_n_n425_ = new_nw_ & new_nv_ & new_n_n19_;
  assign new_n_n417_ = new_ny_ & new_nu_ & new_n_n21_;
  assign new_n_n412_ = new_n_n61_ & new_n_n140_;
  assign new_ng2_ = new_nd0_ & new_n_n131_;
  assign new_n_n399_ = new_nd0_ & new_n_n29_;
  assign new_n_n391_ = new_ns_ & new_nr_ & new_nv_;
  assign new_n_n377_ = new_nw_ & new_nt_ & new_n_n32_;
  assign new_nw2_ = new_nf0_ & new_n_n161_ & new_n_n39_;
  assign new_n_n356_ = new_n_n42_ & new_n_n140_ & new_n_n41_;
  assign new_n_n352_ = new_ns_ & new_ny_;
  assign new_ng3_ = new_n_n143_ & new_n_n46_;
  assign new_n_n340_ = new_n_n129_ & new_n_n63_;
  assign new_n_n331_ = new_n_n48_ & new_n_n124_ & new_n_n47_;
  assign new_n_n325_ = new_n_n52_ & new_n_n121_ & new_n_n50_;
  assign new_n_n315_ = new_ny_ & new_nx_ & new_nw_;
  assign new_n_n307_ = new_n_n64_ & new_nh0_;
  assign new_nc4_ = new_n_n299_ | new_n_n297_ | new_n_n296_ | new_n_n295_ | new_n_n298_ | new_n_n300_;
  assign new_nd4_ = new_nc0_ | new_nd0_;
  assign new_nl4_ = new_nr_ & new_n_n142_ & new_n_n79_;
  assign new_n_n289_ = new_nf0_ & new_ne0_ & new_n_n115_;
  assign new_n_n283_ = new_n_n89_ & new_n_n122_;
  assign new_n_n279_ = new_ne0_ & new_n_n122_ & new_n_n90_;
  assign new_ng5_ = new_nf0_ | new_n_n223_ | new_n_n222_;
  assign new_n_n268_ = new_n_n98_ & new_n_n107_ & new_n_n96_;
  assign new_n_n261_ = new_nq_ & new_n_n105_ & new_n_n104_;
  assign new_n_n252_ = new_n_n116_ & new_nt_;
  assign new_nb6_ = new_n_n122_ | new_n_n121_;
  assign new_n_n242_ = new_nd0_ & new_ne0_;
  assign new_n_n236_ = new_n_n131_ & new_nt_ & new_n_n132_;
  assign new_nl6_ = new_n_n230_ | new_n_n135_;
  assign new_np6_ = new_ns_ & new_nr_ & new_n_n142_;
  assign new_n_n220_ = new_n_n144_ & new_n_n161_;
  assign new_n_n212_ = new_n_n159_ & new_nd_ & new_n_n147_;
  assign new_nb7_ = new_n_n197_ | new_n_n196_ | new_n_n195_;
  assign new_n_n186_ = new_n_n165_ & new_n_n164_ & new_n_n156_;
  assign new_n_n176_ = new_ne_ & new_n_n159_ & new_nh_;
  assign new_n_n171_ = new_nf_ & new_n_n161_;
  assign new_n_n163_ = ~new_ne_;
  assign new_n_n156_ = ~new_nq7_;
  assign new_n_n145_ = ~new_ni0_;
  assign new_n_n138_ = ~new_no6_;
  assign new_n_n127_ = ~new_ng6_;
  assign new_n_n3_ = ~new_nf1_;
  assign new_n_n437_ = new_np_ & new_nv_ & new_nw_;
  assign new_n_n430_ = new_n_n36_ & new_n_n16_;
  assign new_n_n424_ = new_nr_ & new_nv_ & new_n_n19_;
  assign new_na2_ = new_n_n415_ | new_n_n417_ | new_n_n414_ | new_n_n416_;
  assign new_nf2_ = new_n_n406_ | new_n_n405_ | new_n_n404_ | new_n_n403_ | new_n_n410_ | new_n_n408_ | new_n_n407_ | new_n_n409_ | new_n_n411_;
  assign new_n_n403_ = new_n_n36_ & new_n_n24_ & new_n_n23_;
  assign new_n_n398_ = new_n_n28_ & new_nc0_;
  assign new_n_n392_ = new_nx_ & new_nw_ & new_nq_;
  assign new_n_n369_ = new_n_n36_ & new_nc_ & new_n_n34_;
  assign new_ny2_ = new_n_n362_ | new_n_n360_ | new_n_n359_ | new_n_n361_ | new_n_n363_;
  assign new_n_n357_ = new_n_n139_ & new_n_n140_ & new_n_n41_;
  assign new_n_n351_ = new_nx_ & new_nt_;
  assign new_n_n345_ = new_nw_ & new_ns_ & new_n_n45_;
  assign new_n_n339_ = new_n_n131_ & new_n_n61_;
  assign new_n_n332_ = new_n_n140_ & new_n_n124_ & new_n_n47_;
  assign new_n_n324_ = new_n_n62_ & new_n_n51_ & new_n_n50_;
  assign new_n_n316_ = new_nt_ & new_nx_ & new_nw_;
  assign new_n_n306_ = new_n_n64_ & new_n_n65_;
  assign new_nb4_ = new_nr_ & new_nq_ & new_n_n79_;
  assign new_ne4_ = new_n_n143_ | new_n_n139_ | new_n_n140_;
  assign new_nk4_ = new_n_n139_ | new_n_n143_;
  assign new_nq4_ = new_nq_ | new_n_n107_ | new_n_n142_;
  assign new_nu4_ = new_n_n283_ | new_n_n282_ | new_n_n281_;
  assign new_n_n278_ = new_ne0_ & new_n_n91_ & new_n_n90_;
  assign new_nf5_ = new_n_n133_ & new_n_n129_;
  assign new_n_n267_ = new_n_n94_ & new_n_n97_ & new_n_n96_;
  assign new_n_n262_ = new_ne0_ & new_n_n103_ & new_n_n102_;
  assign new_n_n251_ = new_nr_ & new_ns_ & new_n_n116_;
  assign new_ny5_ = new_n_n143_ | new_n_n139_ | new_nm_;
  assign new_nf6_ = new_ng0_ | new_nf0_ | new_n_n127_;
  assign new_nj6_ = new_n_n234_ | new_n_n236_ | new_n_n233_ | new_n_n235_;
  assign new_n_n230_ = new_n_n136_ & new_n_n140_;
  assign new_no6_ = new_n_n141_ | new_n_n143_;
  assign new_n_n219_ = new_n_n144_ & new_nc_;
  assign new_n_n213_ = new_n_n149_ & new_n_n165_ & new_n_n147_;
  assign new_n_n205_ = new_n_n150_ & new_nc_;
  assign new_n_n185_ = new_nd_ & new_n_n164_ & new_n_n156_;
  assign new_n_n177_ = new_nc_ & new_ne_ & new_nh_;
  assign new_n_n170_ = new_ng_ & new_n_n162_;
  assign new_n_n164_ = ~new_nh_;
  assign new_n_n155_ = ~new_ng7_;
  assign new_n_n146_ = ~new_ni_;
  assign new_n_n137_ = ~new_nn6_;
  assign new_n_n128_ = ~new_nh6_;
  assign new_n_n4_ = ~new_ne1_;
  assign new_n_n93_ = ~new_nb5_;
  assign new_n_n82_ = ~new_ng5_;
  assign new_n_n71_ = ~new_na4_;
  assign new_n_n61_ = ~new_nw_;
  assign new_n_n50_ = ~new_no3_;
  assign new_n_n94_ = ~new_ni5_;
  assign new_n_n81_ = ~new_no_;
  assign new_n_n72_ = ~new_nb4_;
  assign new_n_n60_ = ~new_nt3_;
  assign new_n_n51_ = ~new_nn3_;
  assign new_n_n95_ = ~new_nj5_;
  assign new_n_n80_ = ~new_nn_;
  assign new_n_n69_ = ~new_np4_;
  assign new_n_n63_ = ~new_nx_;
  assign new_n_n52_ = ~new_nm3_;
  assign new_n_n96_ = ~new_nn5_;
  assign new_n_n79_ = ~new_nk4_;
  assign new_n_n70_ = ~new_nc4_;
  assign new_n_n62_ = ~new_nv_;
  assign new_n_n53_ = ~new_nr3_;
  assign new_n_n0_ = ~new_nt6_;
  assign new_n_n97_ = ~new_nm5_;
  assign new_n_n43_ = ~new_ni3_;
  assign new_n_n32_ = ~new_ns2_;
  assign new_n_n21_ = ~new_nd2_;
  assign new_n_n10_ = ~new_nk3_;
  assign new_n_n98_ = ~new_nk5_;
  assign new_n_n42_ = ~new_nb3_;
  assign new_n_n33_ = ~new_nu2_;
  assign new_n_n20_ = ~new_ne2_;
  assign new_n_n11_ = ~new_nj3_;
  assign new_n_n41_ = ~new_nd3_;
  assign new_n_n30_ = ~new_nq2_;
  assign new_n_n23_ = ~new_ni2_;
  assign new_n_n12_ = ~new_nw3_;
  assign new_n_n40_ = ~new_na3_;
  assign new_n_n31_ = ~new_nn2_;
  assign new_n_n22_ = ~new_ng2_;
  assign new_n_n13_ = ~new_nh5_;
  assign new_n_n68_ = ~new_nq4_;
  assign new_n_n58_ = ~new_na0_;
  assign new_n_n47_ = ~new_ns3_;
  assign new_n_n36_ = ~new_nw1_;
  assign new_n_n25_ = ~new_nr2_;
  assign new_n_n14_ = ~new_nh1_;
  assign new_n_n67_ = ~new_no4_;
  assign new_n_n59_ = ~new_nz2_;
  assign new_n_n46_ = ~new_ny_;
  assign new_n_n37_ = ~new_nf3_;
  assign new_n_n24_ = ~new_nh2_;
  assign new_n_n15_ = ~new_nj1_;
  assign new_n_n88_ = ~new_nt4_;
  assign new_n_n77_ = ~new_ni4_;
  assign new_n_n45_ = ~new_ng3_;
  assign new_n_n34_ = ~new_nw2_;
  assign new_n_n27_ = ~new_nk2_;
  assign new_n_n16_ = ~new_nu1_;
  assign new_n_n87_ = ~new_nw4_;
  assign new_n_n78_ = ~new_nj4_;
  assign new_n_n44_ = ~new_nh3_;
  assign new_n_n35_ = ~new_nv2_;
  assign new_n_n26_ = ~new_nz1_;
  assign new_n_n17_ = ~new_na2_;
  assign new_n_n89_ = ~new_nc5_;
  assign new_n_n86_ = ~new_nx4_;
  assign new_n_n75_ = ~new_ng4_;
  assign new_n_n64_ = ~new_nz3_;
  assign new_n_n54_ = ~new_nb_;
  assign new_n_n29_ = ~new_nl2_;
  assign new_n_n18_ = ~new_nx1_;
  assign new_n_n90_ = ~new_ny4_;
  assign new_n_n85_ = ~new_ns4_;
  assign new_n_n76_ = ~new_nh4_;
  assign new_nj0_ = ~new_nh0_;
  assign new_n_n55_ = ~new_nz_;
  assign new_n_n28_ = ~new_nm2_;
  assign new_n_n19_ = ~new_ny1_;
  assign new_n_n91_ = ~new_nd4_;
  assign new_n_n84_ = ~new_nv4_;
  assign new_n_n73_ = ~new_nl4_;
  assign new_n_n66_ = ~new_nr4_;
  assign new_n_n56_ = ~new_np3_;
  assign new_n_n49_ = ~new_nu_;
  assign new_n_n38_ = ~new_ne3_;
  assign new_n_n92_ = ~new_nz4_;
  assign new_n_n83_ = ~new_nu4_;
  assign new_n_n74_ = ~new_nf4_;
  assign new_n_n65_ = ~new_ny3_;
  assign new_n_n57_ = ~new_nq3_;
  assign new_n_n48_ = ~new_nc3_;
  assign new_n_n39_ = ~new_ny2_;
endmodule


