// Benchmark "top" written by ABC on Fri Mar 31 12:12:11 2023

module top ( 
    pv47_3_, pv84_15_, pv84_26_, pv116_20_, pv133_10_, pv15_9_, pv15_14_,
    pv47_4_, pv84_16_, pv84_25_, pv116_9_, pv116_21_, pv119_0_, pv15_13_,
    pv47_5_, pv84_13_, pv84_24_, pv15_12_, pv47_6_, pv84_14_, pv84_23_,
    pv15_6_, pv47_7_, pv47_18_, pv47_29_, pv84_6_, pv84_19_, pv116_6_,
    pv116_11_, pv118_0_, pv15_5_, pv47_8_, pv47_17_, pv84_7_, pv84_29_,
    pv116_5_, pv116_10_, pv15_8_, pv47_9_, pv47_27_, pv84_8_, pv84_17_,
    pv84_28_, pv116_8_, pv15_7_, pv47_19_, pv47_28_, pv84_9_, pv84_18_,
    pv84_27_, pv116_7_, pv118_1_, pv47_14_, pv47_25_, pv116_15_, pv116_28_,
    pv47_13_, pv47_26_, pv84_30_, pv116_14_, pv116_29_, pv122_0_, pv47_16_,
    pv47_23_, pv84_31_, pv116_13_, pv116_26_, pv47_15_, pv47_24_,
    pv116_12_, pv116_27_, pv15_11_, pv47_10_, pv47_21_, pv84_11_, pv84_22_,
    pv116_19_, pv116_24_, pv15_10_, pv47_22_, pv47_31_, pv84_12_, pv84_21_,
    pv116_18_, pv116_25_, pv47_12_, pv47_30_, pv84_20_, pv116_17_,
    pv116_22_, pv116_31_, pv47_11_, pv47_20_, pv84_10_, pv116_16_,
    pv116_23_, pv116_30_, pv133_5_, pv52_0_, pv133_4_, pv133_3_, pv133_2_,
    pv133_1_, pv133_0_, pv15_2_, pv84_2_, pv116_2_, pv121_17_, pv15_1_,
    pv84_3_, pv116_1_, pv15_4_, pv84_4_, pv116_4_, pv15_3_, pv84_5_,
    pv116_3_, pv121_16_, pv133_9_, pv47_0_, pv133_8_, pv15_0_, pv47_1_,
    pv48_0_, pv51_0_, pv84_0_, pv116_0_, pv133_7_, pv47_2_, pv49_0_,
    pv50_0_, pv84_1_, pv133_6_,
    pv150_0_, pv197_21_, pv197_20_, pv197_10_, pv197_11_, pv212_9_,
    pv212_8_, pv142_0_, pv197_7_, pv197_6_, pv165_8_, pv197_9_, pv165_9_,
    pv197_8_, pv149_0_, pv197_3_, pv149_1_, pv197_2_, pv149_2_, pv197_5_,
    pv197_4_, pv145_0_, pv165_2_, pv212_14_, pv145_1_, pv165_3_, pv165_10_,
    pv134_0_, pv165_0_, pv197_1_, pv212_12_, pv146_0_, pv165_1_, pv197_0_,
    pv212_13_, pv165_6_, pv165_13_, pv165_7_, pv165_14_, pv165_4_,
    pv165_11_, pv165_5_, pv165_12_, pv142_1_, pv197_16_, pv197_29_,
    pv212_5_, pv142_2_, pv197_17_, pv197_28_, pv212_4_, pv142_3_, pv143_0_,
    pv197_18_, pv197_27_, pv212_7_, pv136_1_, pv142_4_, pv197_19_,
    pv197_26_, pv212_6_, pv214_0_, pv136_0_, pv142_5_, pv197_12_,
    pv197_25_, pv197_30_, pv212_1_, pv212_10_, pv197_13_, pv197_24_,
    pv197_31_, pv212_0_, pv212_11_, pv197_14_, pv197_23_, pv212_3_,
    pv213_0_, pv197_15_, pv197_22_, pv212_2_  );
  input  pv47_3_, pv84_15_, pv84_26_, pv116_20_, pv133_10_, pv15_9_,
    pv15_14_, pv47_4_, pv84_16_, pv84_25_, pv116_9_, pv116_21_, pv119_0_,
    pv15_13_, pv47_5_, pv84_13_, pv84_24_, pv15_12_, pv47_6_, pv84_14_,
    pv84_23_, pv15_6_, pv47_7_, pv47_18_, pv47_29_, pv84_6_, pv84_19_,
    pv116_6_, pv116_11_, pv118_0_, pv15_5_, pv47_8_, pv47_17_, pv84_7_,
    pv84_29_, pv116_5_, pv116_10_, pv15_8_, pv47_9_, pv47_27_, pv84_8_,
    pv84_17_, pv84_28_, pv116_8_, pv15_7_, pv47_19_, pv47_28_, pv84_9_,
    pv84_18_, pv84_27_, pv116_7_, pv118_1_, pv47_14_, pv47_25_, pv116_15_,
    pv116_28_, pv47_13_, pv47_26_, pv84_30_, pv116_14_, pv116_29_,
    pv122_0_, pv47_16_, pv47_23_, pv84_31_, pv116_13_, pv116_26_, pv47_15_,
    pv47_24_, pv116_12_, pv116_27_, pv15_11_, pv47_10_, pv47_21_, pv84_11_,
    pv84_22_, pv116_19_, pv116_24_, pv15_10_, pv47_22_, pv47_31_, pv84_12_,
    pv84_21_, pv116_18_, pv116_25_, pv47_12_, pv47_30_, pv84_20_,
    pv116_17_, pv116_22_, pv116_31_, pv47_11_, pv47_20_, pv84_10_,
    pv116_16_, pv116_23_, pv116_30_, pv133_5_, pv52_0_, pv133_4_, pv133_3_,
    pv133_2_, pv133_1_, pv133_0_, pv15_2_, pv84_2_, pv116_2_, pv121_17_,
    pv15_1_, pv84_3_, pv116_1_, pv15_4_, pv84_4_, pv116_4_, pv15_3_,
    pv84_5_, pv116_3_, pv121_16_, pv133_9_, pv47_0_, pv133_8_, pv15_0_,
    pv47_1_, pv48_0_, pv51_0_, pv84_0_, pv116_0_, pv133_7_, pv47_2_,
    pv49_0_, pv50_0_, pv84_1_, pv133_6_;
  output pv150_0_, pv197_21_, pv197_20_, pv197_10_, pv197_11_, pv212_9_,
    pv212_8_, pv142_0_, pv197_7_, pv197_6_, pv165_8_, pv197_9_, pv165_9_,
    pv197_8_, pv149_0_, pv197_3_, pv149_1_, pv197_2_, pv149_2_, pv197_5_,
    pv197_4_, pv145_0_, pv165_2_, pv212_14_, pv145_1_, pv165_3_, pv165_10_,
    pv134_0_, pv165_0_, pv197_1_, pv212_12_, pv146_0_, pv165_1_, pv197_0_,
    pv212_13_, pv165_6_, pv165_13_, pv165_7_, pv165_14_, pv165_4_,
    pv165_11_, pv165_5_, pv165_12_, pv142_1_, pv197_16_, pv197_29_,
    pv212_5_, pv142_2_, pv197_17_, pv197_28_, pv212_4_, pv142_3_, pv143_0_,
    pv197_18_, pv197_27_, pv212_7_, pv136_1_, pv142_4_, pv197_19_,
    pv197_26_, pv212_6_, pv214_0_, pv136_0_, pv142_5_, pv197_12_,
    pv197_25_, pv197_30_, pv212_1_, pv212_10_, pv197_13_, pv197_24_,
    pv197_31_, pv212_0_, pv212_11_, pv197_14_, pv197_23_, pv212_3_,
    pv213_0_, pv197_15_, pv197_22_, pv212_2_;
  wire new_n_n245_, new_n_n199_, new_n_n210_, new_n_n160_, new_n_n277_,
    new_n_n225_, new_n_n230_, new_n_n246_, new_n_n200_, new_n_n209_,
    new_n_n179_, new_n_n161_, new_n_n155_, new_n_n229_, new_n_n247_,
    new_n_n197_, new_n_n208_, new_n_n228_, new_n_n248_, new_n_n198_,
    new_n_n207_, new_n_n222_, new_n_n249_, new_n_n260_, new_n_n271_,
    new_n_n236_, new_n_n203_, new_n_n183_, new_n_n178_, new_n_n151_,
    new_n_n221_, new_n_n250_, new_n_n259_, new_n_n237_, new_n_n213_,
    new_n_n182_, new_n_n177_, new_n_n224_, new_n_n251_, new_n_n269_,
    new_n_n238_, new_n_n201_, new_n_n212_, new_n_n185_, new_n_n223_,
    new_n_n261_, new_n_n270_, new_n_n239_, new_n_n202_, new_n_n211_,
    new_n_n184_, new_n_n150_, new_n_n256_, new_n_n267_, new_n_n175_,
    new_n_n168_, new_n_n255_, new_n_n268_, new_n_n214_, new_n_n174_,
    new_n_n169_, new_n_n153_, new_n_n258_, new_n_n265_, new_n_n215_,
    new_n_n173_, new_n_n166_, new_n_n257_, new_n_n266_, new_n_n176_,
    new_n_n167_, new_n_n227_, new_n_n252_, new_n_n263_, new_n_n241_,
    new_n_n206_, new_n_n159_, new_n_n164_, new_n_n226_, new_n_n264_,
    new_n_n273_, new_n_n196_, new_n_n205_, new_n_n158_, new_n_n165_,
    new_n_n254_, new_n_n272_, new_n_n204_, new_n_n157_, new_n_n162_,
    new_n_n171_, new_n_n253_, new_n_n262_, new_n_n240_, new_n_n172_,
    new_n_n163_, new_n_n170_, new_n_n278_, new_n_n190_, new_n_n152_,
    new_n_n282_, new_n_n280_, new_n_n281_, new_n_n279_, new_n_n218_,
    new_n_n232_, new_n_n188_, new_n_n154_, new_n_n217_, new_n_n233_,
    new_n_n186_, new_n_n220_, new_n_n234_, new_n_n181_, new_n_n219_,
    new_n_n235_, new_n_n180_, new_n_n156_, new_n_n187_, new_n_n242_,
    new_n_n274_, new_n_n216_, new_n_n243_, new_n_n194_, new_n_n189_,
    new_n_n195_, new_n_n192_, new_n_n275_, new_n_n244_, new_n_n193_,
    new_n_n191_, new_n_n231_, new_n_n276_, new_nv226_, new_nv238_,
    new_n_n57_, new_nv294_, new_n_n46_, new_n_n40_, new_nv328_, new_nv339_,
    new_nv362_, new_nv397_, new_nv408_, new_nv419_, new_n_n29_, new_nv442_,
    new_n_n18_, new_nv464_, new_n_n7_, new_nv498_, new_nv509_, new_nv521_,
    new_nv532_, new_nv543_, new_nv558_, new_n_n147_, new_nv595_,
    new_nv605_, new_nv614_, new_nv630_, new_nv645_, new_nv668_, new_nv680_,
    new_nv698_, new_nv719_, new_nv730_, new_nv738_, new_n_n122_,
    new_nv752_, new_nv763_, new_nv776_, new_nv788_, new_nv801_, new_nv812_,
    new_nv824_, new_nv836_, new_nv847_, new_n_n115_, new_nv874_,
    new_n_n104_, new_nv885_, new_n_n93_, new_nv896_, new_nv907_,
    new_nv918_, new_nv953_, new_nv964_, new_nv977_, new_nv988_, new_nv999_,
    new_nv1011_, new_nv1022_, new_nv1068_, new_nv1079_, new_nv1088_,
    new_n_n76_, new_nv1100_, new_nv1111_, new_nv228_, new_nv237_,
    new_nv284_, new_n_n52_, new_nv306_, new_n_n41_, new_nv329_, new_nv338_,
    new_nv372_, new_nv398_, new_nv407_, new_nv420_, new_nv430_, new_n_n23_,
    new_nv452_, new_n_n12_, new_nv474_, new_nv499_, new_nv508_, new_nv522_,
    new_nv531_, new_nv544_, new_nv555_, new_nv577_, new_nv594_, new_nv613_,
    new_nv616_, new_nv628_, new_nv648_, new_nv665_, new_nv682_, new_nv695_,
    new_nv720_, new_nv729_, new_n_n127_, new_nv743_, new_nv744_,
    new_nv764_, new_nv775_, new_nv789_, new_nv800_, new_nv813_, new_nv823_,
    new_nv837_, new_nv846_, new_nv869_, new_n_n110_, new_nv880_,
    new_n_n99_, new_nv891_, new_n_n88_, new_nv908_, new_nv917_, new_nv943_,
    new_nv965_, new_nv976_, new_nv989_, new_nv998_, new_nv1012_,
    new_nv1021_, new_nv1069_, new_nv1078_, new_n_n81_, new_nv1093_,
    new_nv1101_, new_nv1110_, new_nv223_, new_nv236_, new_n_n58_,
    new_nv292_, new_n_n45_, new_n_n38_, new_nv326_, new_nv337_, new_nv382_,
    new_nv395_, new_nv406_, new_nv422_, new_n_n28_, new_nv440_, new_n_n19_,
    new_nv484_, new_nv496_, new_nv507_, new_nv523_, new_nv534_, new_nv541_,
    new_nv553_, new_nv578_, new_nv604_, new_nv612_, new_n_n137_,
    new_nv669_, new_nv678_, new_nv693_, new_nv721_, new_n_n132_,
    new_nv737_, new_n_n123_, new_nv767_, new_nv778_, new_nv786_,
    new_nv797_, new_nv814_, new_nv826_, new_nv834_, new_nv845_,
    new_n_n114_, new_nv875_, new_n_n105_, new_nv884_, new_n_n92_,
    new_nv897_, new_nv905_, new_nv916_, new_nv944_, new_nv955_, new_nv975_,
    new_nv990_, new_nv1002_, new_nv1009_, new_nv1020_, new_nv1047_,
    new_nv1058_, new_nv1089_, new_n_n75_, new_nv1098_, new_nv1109_,
    new_nv224_, new_n_n65_, new_nv282_, new_n_n53_, new_nv308_, new_n_n39_,
    new_nv327_, new_nv336_, new_nv394_, new_nv396_, new_nv405_, new_n_n33_,
    new_nv432_, new_n_n24_, new_nv450_, new_n_n2_, new_nv495_, new_nv497_,
    new_nv524_, new_nv533_, new_nv542_, new_nv551_, new_nv596_,
    new_n_n144_, new_nv611_, new_nv651_, new_n_n136_, new_nv679_,
    new_nv692_, new_nv722_, new_nv733_, new_n_n128_, new_nv742_,
    new_nv768_, new_nv777_, new_nv787_, new_nv796_, new_nv816_, new_nv825_,
    new_nv835_, new_nv844_, new_nv870_, new_n_n109_, new_nv879_,
    new_n_n100_, new_nv892_, new_n_n87_, new_nv906_, new_nv915_,
    new_nv945_, new_nv954_, new_nv963_, new_nv991_, new_nv1001_,
    new_nv1010_, new_nv1019_, new_nv1048_, new_nv1057_, new_n_n80_,
    new_nv1094_, new_n_n71_, new_nv1108_, new_nv219_, new_n_n66_,
    new_n_n55_, new_nv298_, new_n_n48_, new_nv312_, new_nv324_, new_nv335_,
    new_nv401_, new_nv412_, new_nv415_, new_n_n31_, new_nv438_, new_n_n20_,
    new_nv502_, new_nv513_, new_nv528_, new_nv539_, new_nv550_, new_nv619_,
    new_n_n139_, new_nv674_, new_nv691_, new_n_n120_, new_nv756_,
    new_nv795_, new_nv817_, new_nv851_, new_nv862_, new_n_n91_, new_nv900_,
    new_nv922_, new_nv935_, new_nv992_, new_nv1004_, new_nv1015_,
    new_nv1026_, new_nv1038_, new_nv1090_, new_n_n74_, new_nv1104_,
    new_nv1117_, new_nv582_, new_nv222_, new_n_n67_, new_nv288_,
    new_n_n50_, new_nv302_, new_n_n43_, new_nv325_, new_nv334_, new_nv402_,
    new_nv411_, new_nv416_, new_nv426_, new_n_n25_, new_nv448_, new_nv503_,
    new_nv512_, new_nv517_, new_nv540_, new_nv549_, new_nv620_, new_nv636_,
    new_nv675_, new_nv689_, new_nv746_, new_nv755_, new_nv785_, new_nv827_,
    new_nv852_, new_nv861_, new_nv893_, new_n_n86_, new_nv923_, new_nv934_,
    new_nv993_, new_nv1003_, new_nv1025_, new_nv1027_, new_nv1037_,
    new_n_n79_, new_nv1095_, new_nv1105_, new_nv1114_, new_n_n68_,
    new_n_n56_, new_nv296_, new_n_n47_, new_nv314_, new_n_n35_, new_nv333_,
    new_nv399_, new_nv410_, new_nv417_, new_n_n30_, new_nv436_, new_n_n21_,
    new_nv500_, new_nv511_, new_nv518_, new_nv530_, new_nv548_, new_nv617_,
    new_nv633_, new_nv642_, new_nv664_, new_n_n121_, new_nv754_,
    new_nv774_, new_nv838_, new_nv849_, new_nv860_, new_nv909_, new_nv920_,
    new_nv931_, new_nv994_, new_nv1013_, new_nv1024_, new_nv1091_,
    new_n_n73_, new_nv1102_, new_nv1113_, new_nv215_, new_nv231_,
    new_nv286_, new_n_n51_, new_nv304_, new_n_n42_, new_n_n34_, new_nv332_,
    new_nv400_, new_nv409_, new_nv418_, new_nv428_, new_n_n26_, new_nv446_,
    new_nv501_, new_nv510_, new_nv520_, new_nv529_, new_nv538_, new_nv618_,
    new_nv632_, new_nv643_, new_nv663_, new_nv745_, new_nv753_, new_nv762_,
    new_nv848_, new_nv850_, new_nv859_, new_nv910_, new_nv919_, new_nv921_,
    new_nv1005_, new_nv1014_, new_nv1023_, new_n_n78_, new_nv1096_,
    new_nv1103_, new_nv1112_, new_nv241_, new_nv252_, new_nv263_,
    new_n_n61_, new_nv342_, new_nv365_, new_nv376_, new_nv389_, new_nv456_,
    new_n_n11_, new_nv478_, new_nv490_, new_nv506_, new_nv581_, new_nv598_,
    new_n_n142_, new_nv626_, new_nv640_, new_nv734_, new_n_n126_,
    new_n_n118_, new_nv760_, new_nv773_, new_nv839_, new_nv855_,
    new_nv867_, new_n_n111_, new_nv878_, new_nv926_, new_nv939_,
    new_nv950_, new_nv961_, new_nv974_, new_nv1030_, new_nv1042_,
    new_nv1053_, new_nv1064_, new_nv1076_, new_n_n83_, new_nv559_,
    new_nv242_, new_nv251_, new_nv264_, new_nv274_, new_nv343_, new_nv364_,
    new_nv377_, new_nv386_, new_n_n16_, new_nv466_, new_n_n5_, new_nv489_,
    new_nv516_, new_nv566_, new_nv599_, new_nv606_, new_n_n140_,
    new_nv639_, new_n_n131_, new_nv739_, new_nv750_, new_nv759_,
    new_nv784_, new_nv828_, new_nv856_, new_n_n117_, new_nv873_,
    new_n_n106_, new_nv927_, new_nv938_, new_nv951_, new_nv960_,
    new_nv984_, new_nv1031_, new_nv1041_, new_nv1054_, new_nv1063_,
    new_nv1077_, new_nv1086_, new_nv562_, new_nv243_, new_nv254_,
    new_nv261_, new_n_n62_, new_n_n54_, new_nv356_, new_nv367_, new_nv374_,
    new_nv385_, new_nv403_, new_nv414_, new_nv458_, new_n_n10_, new_nv476_,
    new_nv488_, new_nv504_, new_nv515_, new_nv568_, new_nv585_,
    new_n_n143_, new_nv621_, new_n_n138_, new_nv709_, new_nv724_,
    new_n_n119_, new_nv758_, new_nv794_, new_nv818_, new_nv853_,
    new_nv866_, new_n_n101_, new_nv888_, new_nv924_, new_nv937_,
    new_nv952_, new_nv972_, new_nv983_, new_nv1028_, new_nv1040_,
    new_nv1055_, new_nv1067_, new_nv1074_, new_n_n84_, new_nv572_,
    new_nv244_, new_nv253_, new_nv262_, new_nv272_, new_n_n49_, new_nv357_,
    new_nv366_, new_nv375_, new_nv384_, new_nv404_, new_nv413_, new_n_n15_,
    new_nv468_, new_n_n6_, new_nv487_, new_nv505_, new_nv514_, new_nv570_,
    new_nv584_, new_nv597_, new_nv623_, new_nv637_, new_nv712_, new_nv723_,
    new_nv747_, new_nv757_, new_nv806_, new_nv807_, new_nv854_, new_nv863_,
    new_nv883_, new_n_n96_, new_nv925_, new_nv936_, new_nv962_, new_nv973_,
    new_nv982_, new_nv1029_, new_nv1039_, new_nv1056_, new_nv1065_,
    new_nv1075_, new_nv1085_, new_nv576_, new_nv245_, new_nv256_,
    new_nv268_, new_n_n59_, new_n_n44_, new_nv358_, new_nv369_, new_nv380_,
    new_nv393_, new_nv424_, new_n_n27_, new_nv460_, new_n_n9_, new_nv482_,
    new_nv494_, new_nv525_, new_nv536_, new_nv547_, new_nv571_, new_nv589_,
    new_nv603_, new_nv610_, new_nv654_, new_nv670_, new_nv687_, new_nv707_,
    new_nv714_, new_nv726_, new_nv736_, new_n_n124_, new_nv769_,
    new_nv780_, new_nv792_, new_nv805_, new_nv808_, new_nv820_, new_nv832_,
    new_nv843_, new_n_n113_, new_nv876_, new_n_n102_, new_nv887_,
    new_n_n95_, new_nv894_, new_nv903_, new_nv914_, new_nv930_, new_nv946_,
    new_nv957_, new_nv970_, new_nv981_, new_nv995_, new_nv1007_,
    new_nv1018_, new_nv1035_, new_nv1046_, new_nv1049_, new_nv1060_,
    new_nv1072_, new_n_n85_, new_nv1097_, new_nv1107_, new_nv486_,
    new_nv246_, new_nv255_, new_n_n64_, new_nv278_, new_n_n37_, new_nv359_,
    new_nv368_, new_nv381_, new_nv392_, new_n_n32_, new_nv434_, new_n_n14_,
    new_nv470_, new_n_n3_, new_nv493_, new_nv526_, new_nv535_, new_nv564_,
    new_nv574_, new_nv588_, new_n_n145_, new_nv609_, new_nv656_,
    new_n_n135_, new_nv688_, new_nv704_, new_nv716_, new_nv725_,
    new_n_n129_, new_nv741_, new_nv770_, new_nv779_, new_nv793_,
    new_nv804_, new_nv809_, new_nv819_, new_nv833_, new_nv842_, new_nv871_,
    new_n_n108_, new_nv882_, new_n_n97_, new_nv889_, new_n_n90_,
    new_nv904_, new_nv913_, new_nv942_, new_nv947_, new_nv956_, new_nv971_,
    new_nv980_, new_nv985_, new_nv1008_, new_nv1017_, new_nv1036_,
    new_nv1045_, new_nv1050_, new_nv1059_, new_nv1073_, new_nv1084_,
    new_n_n72_, new_nv1106_, new_nv519_, new_nv247_, new_nv258_,
    new_nv265_, new_n_n60_, new_nv330_, new_nv360_, new_nv371_, new_nv378_,
    new_nv391_, new_nv444_, new_n_n17_, new_nv462_, new_n_n8_, new_nv480_,
    new_nv492_, new_nv527_, new_nv545_, new_nv561_, new_n_n148_,
    new_nv592_, new_nv602_, new_n_n141_, new_nv659_, new_nv673_,
    new_nv683_, new_nv701_, new_nv717_, new_nv728_, new_nv735_,
    new_n_n125_, new_nv751_, new_nv771_, new_nv783_, new_nv790_,
    new_nv803_, new_nv810_, new_nv822_, new_nv829_, new_nv841_, new_nv857_,
    new_nv868_, new_n_n112_, new_nv877_, new_n_n103_, new_nv886_,
    new_n_n94_, new_nv895_, new_nv901_, new_nv912_, new_nv928_, new_nv941_,
    new_nv948_, new_nv959_, new_nv968_, new_nv979_, new_nv986_, new_nv997_,
    new_nv1016_, new_nv1032_, new_nv1044_, new_nv1051_, new_nv1062_,
    new_nv1070_, new_nv1081_, new_nv1087_, new_n_n77_, new_nv552_,
    new_nv248_, new_nv257_, new_nv266_, new_nv276_, new_nv340_, new_nv361_,
    new_nv370_, new_nv379_, new_nv390_, new_n_n22_, new_nv454_, new_n_n13_,
    new_nv472_, new_n_n4_, new_nv491_, new_nv537_, new_nv546_, new_n_n149_,
    new_nv575_, new_nv591_, new_n_n146_, new_nv607_, new_nv661_,
    new_n_n134_, new_nv684_, new_n_n133_, new_nv718_, new_nv727_,
    new_n_n130_, new_nv740_, new_nv761_, new_nv772_, new_nv781_,
    new_nv791_, new_nv802_, new_nv811_, new_nv821_, new_nv830_, new_nv840_,
    new_nv858_, new_n_n116_, new_nv872_, new_n_n107_, new_nv881_,
    new_n_n98_, new_nv890_, new_n_n89_, new_nv902_, new_nv911_, new_nv929_,
    new_nv940_, new_nv949_, new_nv958_, new_nv969_, new_nv978_, new_nv987_,
    new_nv996_, new_nv1006_, new_nv1034_, new_nv1043_, new_nv1052_,
    new_nv1061_, new_nv1071_, new_nv1080_, new_n_n82_, new_nv1092_,
    new_nv556_, new_nv1124_, new_n_n70_, new_nv560_, new_nv749_,
    new_nv1139_, new_nv1123_, new_nv1141_, new_nv557_, new_nv799_,
    new_nv1134_, new_nv1122_, new_nv1144_, new_nv573_, new_nv706_,
    new_nv1116_, new_nv1121_, new_nv1147_, new_nv569_, new_nv732_,
    new_nv1083_, new_nv421_, new_nv259_, new_n_n63_, new_nv383_,
    new_nv1120_, new_nv1310_, new_nv1155_, new_nv864_, new_nv586_,
    new_nv260_, new_nv270_, new_nv373_, new_nv1119_, new_nv1309_,
    new_nv1263_, new_nv699_, new_nv590_, new_nv239_, new_nv250_,
    new_nv363_, new_nv1302_, new_nv1140_, new_nv932_, new_nv600_,
    new_nv240_, new_nv249_, new_nv341_, new_nv1300_, new_nv1152_,
    new_nv898_, new_nv624_, new_nv230_, new_nv331_, new_nv587_, new_nv865_,
    new_nv1150_, new_nv1288_, new_nv1000_, new_nv627_, new_nv229_,
    new_n_n36_, new_nv622_, new_nv831_, new_nv1153_, new_nv1289_,
    new_nv966_, new_nv646_, new_nv310_, new_nv1129_, new_nv1151_,
    new_nv1316_, new_nv1276_, new_nv1099_, new_nv649_, new_nv300_,
    new_nv1130_, new_nv1149_, new_nv1315_, new_nv1287_, new_nv1082_,
    new_nv652_, new_nv290_, new_nv1128_, new_nv1131_, new_n_n69_,
    new_nv694_, new_nv1066_, new_nv1136_, new_nv660_, new_nv280_,
    new_nv1127_, new_nv1132_, new_nv1154_, new_nv697_, new_nv967_,
    new_nv1118_, new_nv696_, new_nv1126_, new_nv1133_, new_nv554_,
    new_nv631_, new_nv933_, new_nv1143_, new_nv1295_, new_nv1125_,
    new_nv1135_, new_nv1156_, new_nv644_, new_nv899_, new_nv1146_,
    new_nv1299_;
  assign new_n_n245_ = pv47_3_;
  assign new_n_n199_ = pv84_15_;
  assign new_n_n210_ = pv84_26_;
  assign new_n_n160_ = pv116_20_;
  assign new_n_n277_ = pv133_10_;
  assign pv150_0_ = new_n_n133_;
  assign pv197_21_ = new_n_n107_;
  assign new_n_n225_ = pv15_9_;
  assign new_n_n230_ = pv15_14_;
  assign new_n_n246_ = pv47_4_;
  assign new_n_n200_ = pv84_16_;
  assign new_n_n209_ = pv84_25_;
  assign new_n_n179_ = pv116_9_;
  assign new_n_n161_ = pv116_21_;
  assign new_n_n155_ = pv119_0_;
  assign pv197_20_ = new_n_n106_;
  assign new_n_n229_ = pv15_13_;
  assign new_n_n247_ = pv47_5_;
  assign new_n_n197_ = pv84_13_;
  assign new_n_n208_ = pv84_24_;
  assign pv197_10_ = new_n_n96_;
  assign new_n_n228_ = pv15_12_;
  assign new_n_n248_ = pv47_6_;
  assign new_n_n198_ = pv84_14_;
  assign new_n_n207_ = pv84_23_;
  assign pv197_11_ = new_n_n97_;
  assign new_n_n222_ = pv15_6_;
  assign new_n_n249_ = pv47_7_;
  assign new_n_n260_ = pv47_18_;
  assign new_n_n271_ = pv47_29_;
  assign new_n_n236_ = pv84_6_;
  assign new_n_n203_ = pv84_19_;
  assign new_n_n183_ = pv116_6_;
  assign new_n_n178_ = pv116_11_;
  assign new_n_n151_ = pv118_0_;
  assign pv212_9_ = new_n_n80_;
  assign new_n_n221_ = pv15_5_;
  assign new_n_n250_ = pv47_8_;
  assign new_n_n259_ = pv47_17_;
  assign new_n_n237_ = pv84_7_;
  assign new_n_n213_ = pv84_29_;
  assign new_n_n182_ = pv116_5_;
  assign new_n_n177_ = pv116_10_;
  assign pv212_8_ = new_n_n79_;
  assign new_n_n224_ = pv15_8_;
  assign new_n_n251_ = pv47_9_;
  assign new_n_n269_ = pv47_27_;
  assign new_n_n238_ = pv84_8_;
  assign new_n_n201_ = pv84_17_;
  assign new_n_n212_ = pv84_28_;
  assign new_n_n185_ = pv116_8_;
  assign new_n_n223_ = pv15_7_;
  assign new_n_n261_ = pv47_19_;
  assign new_n_n270_ = pv47_28_;
  assign new_n_n239_ = pv84_9_;
  assign new_n_n202_ = pv84_18_;
  assign new_n_n211_ = pv84_27_;
  assign new_n_n184_ = pv116_7_;
  assign new_n_n150_ = pv118_1_;
  assign pv142_0_ = new_n_n141_;
  assign new_n_n256_ = pv47_14_;
  assign new_n_n267_ = pv47_25_;
  assign new_n_n175_ = pv116_15_;
  assign new_n_n168_ = pv116_28_;
  assign pv197_7_ = new_n_n93_;
  assign new_n_n255_ = pv47_13_;
  assign new_n_n268_ = pv47_26_;
  assign new_n_n214_ = pv84_30_;
  assign new_n_n174_ = pv116_14_;
  assign new_n_n169_ = pv116_29_;
  assign new_n_n153_ = pv122_0_;
  assign pv197_6_ = new_n_n92_;
  assign new_n_n258_ = pv47_16_;
  assign new_n_n265_ = pv47_23_;
  assign new_n_n215_ = pv84_31_;
  assign new_n_n173_ = pv116_13_;
  assign new_n_n166_ = pv116_26_;
  assign pv165_8_ = new_n_n126_;
  assign pv197_9_ = new_n_n95_;
  assign new_n_n257_ = pv47_15_;
  assign new_n_n266_ = pv47_24_;
  assign new_n_n176_ = pv116_12_;
  assign new_n_n167_ = pv116_27_;
  assign pv165_9_ = new_n_n127_;
  assign pv197_8_ = new_n_n94_;
  assign new_n_n227_ = pv15_11_;
  assign new_n_n252_ = pv47_10_;
  assign new_n_n263_ = pv47_21_;
  assign new_n_n241_ = pv84_11_;
  assign new_n_n206_ = pv84_22_;
  assign new_n_n159_ = pv116_19_;
  assign new_n_n164_ = pv116_24_;
  assign pv149_0_ = new_n_n134_;
  assign pv197_3_ = new_n_n89_;
  assign new_n_n226_ = pv15_10_;
  assign new_n_n264_ = pv47_22_;
  assign new_n_n273_ = pv47_31_;
  assign new_n_n196_ = pv84_12_;
  assign new_n_n205_ = pv84_21_;
  assign new_n_n158_ = pv116_18_;
  assign new_n_n165_ = pv116_25_;
  assign pv149_1_ = new_n_n135_;
  assign pv197_2_ = new_n_n88_;
  assign new_n_n254_ = pv47_12_;
  assign new_n_n272_ = pv47_30_;
  assign new_n_n204_ = pv84_20_;
  assign new_n_n157_ = pv116_17_;
  assign new_n_n162_ = pv116_22_;
  assign new_n_n171_ = pv116_31_;
  assign pv149_2_ = new_n_n136_;
  assign pv197_5_ = new_n_n91_;
  assign new_n_n253_ = pv47_11_;
  assign new_n_n262_ = pv47_20_;
  assign new_n_n240_ = pv84_10_;
  assign new_n_n172_ = pv116_16_;
  assign new_n_n163_ = pv116_23_;
  assign new_n_n170_ = pv116_30_;
  assign pv197_4_ = new_n_n90_;
  assign new_n_n278_ = pv133_5_;
  assign pv145_0_ = new_n_n138_;
  assign pv165_2_ = new_n_n120_;
  assign pv212_14_ = new_n_n85_;
  assign new_n_n190_ = pv52_0_;
  assign new_n_n152_ = pv133_4_;
  assign pv145_1_ = new_n_n139_;
  assign pv165_3_ = new_n_n121_;
  assign pv165_10_ = new_n_n128_;
  assign new_n_n282_ = pv133_3_;
  assign pv134_0_ = new_n_n149_;
  assign pv165_0_ = new_n_n118_;
  assign pv197_1_ = new_n_n87_;
  assign pv212_12_ = new_n_n83_;
  assign new_n_n280_ = pv133_2_;
  assign pv146_0_ = new_n_n137_;
  assign pv165_1_ = new_n_n119_;
  assign pv197_0_ = new_n_n86_;
  assign pv212_13_ = new_n_n84_;
  assign new_n_n281_ = pv133_1_;
  assign pv165_6_ = new_n_n124_;
  assign pv165_13_ = new_n_n131_;
  assign new_n_n279_ = pv133_0_;
  assign pv165_7_ = new_n_n125_;
  assign pv165_14_ = new_n_n132_;
  assign pv165_4_ = new_n_n122_;
  assign pv165_11_ = new_n_n129_;
  assign pv165_5_ = new_n_n123_;
  assign pv165_12_ = new_n_n130_;
  assign new_n_n218_ = pv15_2_;
  assign new_n_n232_ = pv84_2_;
  assign new_n_n188_ = pv116_2_;
  assign new_n_n154_ = pv121_17_;
  assign pv142_1_ = new_n_n142_;
  assign pv197_16_ = new_n_n102_;
  assign pv197_29_ = new_n_n115_;
  assign pv212_5_ = new_n_n76_;
  assign new_n_n217_ = pv15_1_;
  assign new_n_n233_ = pv84_3_;
  assign new_n_n186_ = pv116_1_;
  assign pv142_2_ = new_n_n143_;
  assign pv197_17_ = new_n_n103_;
  assign pv197_28_ = new_n_n114_;
  assign pv212_4_ = new_n_n75_;
  assign new_n_n220_ = pv15_4_;
  assign new_n_n234_ = pv84_4_;
  assign new_n_n181_ = pv116_4_;
  assign pv142_3_ = new_n_n144_;
  assign pv143_0_ = new_n_n140_;
  assign pv197_18_ = new_n_n104_;
  assign pv197_27_ = new_n_n113_;
  assign pv212_7_ = new_n_n78_;
  assign new_n_n219_ = pv15_3_;
  assign new_n_n235_ = pv84_5_;
  assign new_n_n180_ = pv116_3_;
  assign new_n_n156_ = pv121_16_;
  assign pv136_1_ = new_n_n148_;
  assign pv142_4_ = new_n_n145_;
  assign pv197_19_ = new_n_n105_;
  assign pv197_26_ = new_n_n112_;
  assign pv212_6_ = new_n_n77_;
  assign pv214_0_ = new_n_n69_;
  assign new_n_n187_ = pv133_9_;
  assign pv136_0_ = new_n_n147_;
  assign pv142_5_ = new_n_n146_;
  assign pv197_12_ = new_n_n98_;
  assign pv197_25_ = new_n_n111_;
  assign pv197_30_ = new_n_n116_;
  assign pv212_1_ = new_n_n72_;
  assign pv212_10_ = new_n_n81_;
  assign new_n_n242_ = pv47_0_;
  assign new_n_n274_ = pv133_8_;
  assign pv197_13_ = new_n_n99_;
  assign pv197_24_ = new_n_n110_;
  assign pv197_31_ = new_n_n117_;
  assign pv212_0_ = new_n_n71_;
  assign pv212_11_ = new_n_n82_;
  assign new_n_n216_ = pv15_0_;
  assign new_n_n243_ = pv47_1_;
  assign new_n_n194_ = pv48_0_;
  assign new_n_n189_ = pv51_0_;
  assign new_n_n195_ = pv84_0_;
  assign new_n_n192_ = pv116_0_;
  assign new_n_n275_ = pv133_7_;
  assign pv197_14_ = new_n_n100_;
  assign pv197_23_ = new_n_n109_;
  assign pv212_3_ = new_n_n74_;
  assign pv213_0_ = new_n_n70_;
  assign new_n_n244_ = pv47_2_;
  assign new_n_n193_ = pv49_0_;
  assign new_n_n191_ = pv50_0_;
  assign new_n_n231_ = pv84_1_;
  assign new_n_n276_ = pv133_6_;
  assign pv197_15_ = new_n_n101_;
  assign pv197_22_ = new_n_n108_;
  assign pv212_2_ = new_n_n73_;
  assign new_nv226_ = new_nv1316_ & new_n_n281_ & new_nv1263_ & new_n_n280_;
  assign new_nv238_ = new_n_n271_ & new_n_n68_;
  assign new_n_n57_ = new_nv331_ | new_nv553_ | new_nv363_ | new_nv282_ | new_nv243_;
  assign new_nv294_ = new_n_n252_ & new_n_n67_ & new_nv421_;
  assign new_n_n46_ = new_nv342_ | new_nv553_ | new_nv374_ | new_nv304_ | new_nv254_;
  assign new_n_n40_ = new_nv260_ | new_nv500_ | new_nv553_ | new_nv380_;
  assign new_nv328_ = new_n_n258_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv339_ = new_n_n247_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv362_ = new_n_n252_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv397_ = new_n_n207_ & new_n_n68_;
  assign new_nv408_ = new_n_n196_ & new_n_n68_;
  assign new_nv419_ = new_n_n231_ & new_n_n68_;
  assign new_n_n29_ = new_nv491_ | new_nv553_ | new_nv524_ | new_nv430_ | new_nv393_;
  assign new_nv442_ = new_n_n197_ & new_n_n67_ & new_nv421_;
  assign new_n_n18_ = new_nv502_ | new_nv553_ | new_nv535_ | new_nv452_ | new_nv404_;
  assign new_nv464_ = new_n_n232_ & new_n_n67_ & new_nv421_;
  assign new_n_n7_ = new_nv513_ | new_nv553_ | new_nv546_ | new_nv474_ | new_nv415_;
  assign new_nv498_ = new_n_n239_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv509_ = new_n_n272_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv521_ = new_n_n199_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv532_ = new_n_n234_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv543_ = new_n_n267_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv558_ = new_n_n194_ & new_nv557_ & new_nv556_;
  assign new_n_n147_ = new_nv581_ | new_nv578_ | new_nv589_ | new_nv585_ | new_nv571_ | new_nv592_ | new_nv575_;
  assign new_nv595_ = new_n_n40_ & new_nv631_;
  assign new_nv605_ = new_n_n38_ & new_nv706_ & new_nv600_;
  assign new_nv614_ = new_n_n36_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_nv630_ = new_nv1316_ & new_n_n179_ & new_nv624_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_nv645_ = new_n_n45_ & new_nv644_;
  assign new_nv668_ = new_n_n48_ & new_nv732_ & new_nv699_;
  assign new_nv680_ = new_n_n46_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv698_ = new_n_n49_ & new_nv697_ & new_nv696_;
  assign new_nv719_ = new_n_n61_ & new_nv697_;
  assign new_nv730_ = new_n_n50_ & new_nv697_;
  assign new_nv738_ = new_n_n59_ & new_nv732_ & new_nv699_;
  assign new_n_n122_ = new_nv777_ | new_nv760_ | new_nv810_ | new_nv793_ | new_nv726_ | new_nv826_ | new_nv743_;
  assign new_nv752_ = new_n_n62_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv763_ = new_n_n51_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv776_ = new_n_n55_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv788_ = new_n_n277_ & new_n_n59_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv801_ = new_nv799_ & new_nv627_ & new_n_n170_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv812_ = new_nv799_ & new_nv627_ & new_n_n159_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv824_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n207_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv836_ = new_n_n29_ & new_nv831_;
  assign new_nv847_ = new_n_n18_ & new_nv831_;
  assign new_n_n115_ = new_nv936_ | new_nv902_ | new_nv1003_ | new_nv970_ | new_nv834_ | new_nv1036_ | new_nv868_;
  assign new_nv874_ = new_n_n25_ & new_nv865_ & new_nv864_;
  assign new_n_n104_ = new_nv947_ | new_nv913_ | new_nv1014_ | new_nv981_ | new_nv845_ | new_nv1047_ | new_nv879_;
  assign new_nv885_ = new_n_n14_ & new_nv865_ & new_nv864_;
  assign new_n_n93_ = new_nv958_ | new_nv924_ | new_nv1025_ | new_nv992_ | new_nv856_ | new_nv1058_ | new_nv890_;
  assign new_nv896_ = new_n_n3_ & new_nv865_ & new_nv864_;
  assign new_nv907_ = new_n_n26_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv918_ = new_n_n15_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv953_ = new_n_n14_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv964_ = new_n_n3_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv977_ = new_nv967_ & new_n_n24_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv988_ = new_nv967_ & new_n_n13_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv999_ = new_nv967_ & new_n_n2_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1011_ = new_n_n277_ & new_nv966_ & new_n_n23_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1022_ = new_n_n277_ & new_nv966_ & new_n_n12_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1068_ = new_n_n214_ & new_nv1066_;
  assign new_nv1079_ = new_n_n203_ & new_nv1066_;
  assign new_nv1088_ = new_n_n211_ & new_nv1083_ & new_nv1082_;
  assign new_n_n76_ = new_nv1109_ | new_nv1128_ | new_nv1117_ | new_nv1093_ | new_nv1076_;
  assign new_nv1100_ = new_n_n215_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv1111_ = new_n_n204_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv228_ = new_nv1289_ & new_nv1316_ & new_nv1309_ & new_nv1288_ & new_n_n279_ & new_n_n280_;
  assign new_nv237_ = new_n_n272_ & new_n_n68_;
  assign new_nv284_ = new_n_n257_ & new_n_n67_ & new_nv421_;
  assign new_n_n52_ = new_nv336_ | new_nv553_ | new_nv368_ | new_nv292_ | new_nv248_;
  assign new_nv306_ = new_n_n246_ & new_n_n67_ & new_nv421_;
  assign new_n_n41_ = new_nv499_ | new_nv553_ | new_nv379_ | new_nv314_ | new_nv259_;
  assign new_nv329_ = new_n_n257_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv338_ = new_n_n248_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv372_ = new_n_n230_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv398_ = new_n_n206_ & new_n_n68_;
  assign new_nv407_ = new_n_n197_ & new_n_n68_;
  assign new_nv420_ = new_n_n195_ & new_n_n68_;
  assign new_nv430_ = new_n_n203_ & new_n_n67_ & new_nv421_;
  assign new_n_n23_ = new_nv497_ | new_nv553_ | new_nv530_ | new_nv442_ | new_nv399_;
  assign new_nv452_ = new_n_n238_ & new_n_n67_ & new_nv421_;
  assign new_n_n12_ = new_nv508_ | new_nv553_ | new_nv541_ | new_nv464_ | new_nv410_;
  assign new_nv474_ = new_n_n271_ & new_n_n67_ & new_nv421_;
  assign new_nv499_ = new_n_n238_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv508_ = new_n_n273_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv522_ = new_n_n198_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv531_ = new_n_n235_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv544_ = new_n_n266_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv555_ = new_n_n194_ & new_nv554_;
  assign new_nv577_ = new_n_n35_ & new_nv572_ & new_n_n277_ & new_nv576_;
  assign new_nv594_ = new_n_n41_ & new_nv631_;
  assign new_nv613_ = new_n_n37_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_nv616_ = new_nv1316_ & new_n_n185_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_nv628_ = new_n_n42_ & new_nv624_ & new_n_n277_ & new_nv627_;
  assign new_nv648_ = new_n_n45_ & new_nv732_ & new_nv646_;
  assign new_nv665_ = new_n_n46_ & new_nv697_;
  assign new_nv682_ = new_n_n277_ & new_n_n48_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv695_ = new_n_n49_ & new_nv694_;
  assign new_nv720_ = new_n_n60_ & new_nv697_;
  assign new_nv729_ = new_n_n51_ & new_nv697_;
  assign new_n_n127_ = new_nv772_ | new_nv755_ | new_nv805_ | new_nv788_ | new_nv721_ | new_nv821_ | new_nv738_;
  assign new_nv743_ = new_n_n54_ & new_nv732_ & new_nv699_;
  assign new_nv744_ = new_n_n53_ & new_nv732_ & new_nv699_;
  assign new_nv764_ = new_n_n50_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv775_ = new_n_n56_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv789_ = new_n_n277_ & new_n_n58_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv800_ = new_nv799_ & new_nv627_ & new_n_n171_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv813_ = new_nv799_ & new_nv627_ & new_n_n158_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv823_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n208_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv837_ = new_n_n28_ & new_nv831_;
  assign new_nv846_ = new_n_n19_ & new_nv831_;
  assign new_nv869_ = new_n_n30_ & new_nv865_ & new_nv864_;
  assign new_n_n110_ = new_nv941_ | new_nv907_ | new_nv1008_ | new_nv975_ | new_nv839_ | new_nv1041_ | new_nv873_;
  assign new_nv880_ = new_n_n19_ & new_nv865_ & new_nv864_;
  assign new_n_n99_ = new_nv952_ | new_nv918_ | new_nv1019_ | new_nv986_ | new_nv850_ | new_nv1052_ | new_nv884_;
  assign new_nv891_ = new_n_n8_ & new_nv865_ & new_nv864_;
  assign new_n_n88_ = new_nv963_ | new_nv929_ | new_nv1030_ | new_nv997_ | new_nv861_ | new_nv1063_ | new_nv895_;
  assign new_nv908_ = new_n_n25_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv917_ = new_n_n16_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv943_ = new_n_n24_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv965_ = new_n_n2_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv976_ = new_nv967_ & new_n_n25_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv989_ = new_nv967_ & new_n_n12_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv998_ = new_nv967_ & new_n_n3_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1012_ = new_n_n277_ & new_nv966_ & new_n_n22_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1021_ = new_n_n277_ & new_nv966_ & new_n_n13_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1069_ = new_n_n213_ & new_nv1066_;
  assign new_nv1078_ = new_n_n204_ & new_nv1066_;
  assign new_n_n81_ = new_nv1104_ | new_nv1123_ | new_nv1117_ | new_nv1088_ | new_nv1071_;
  assign new_nv1093_ = new_n_n206_ & new_nv1083_ & new_nv1082_;
  assign new_nv1101_ = new_n_n214_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv1110_ = new_n_n205_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv223_ = new_nv1316_ & new_nv1276_ & new_n_n275_;
  assign new_nv236_ = new_n_n273_ & new_n_n68_;
  assign new_n_n58_ = new_nv330_ | new_nv553_ | new_nv362_ | new_nv280_ | new_nv242_;
  assign new_nv292_ = new_n_n253_ & new_n_n67_ & new_nv421_;
  assign new_n_n45_ = new_nv343_ | new_nv553_ | new_nv375_ | new_nv306_ | new_nv255_;
  assign new_n_n38_ = new_nv262_ | new_nv502_ | new_nv553_ | new_nv382_;
  assign new_nv326_ = new_n_n260_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv337_ = new_n_n249_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv382_ = new_n_n220_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv395_ = new_n_n209_ & new_n_n68_;
  assign new_nv406_ = new_n_n198_ & new_n_n68_;
  assign new_nv422_ = new_n_n207_ & new_n_n67_ & new_nv421_;
  assign new_n_n28_ = new_nv492_ | new_nv553_ | new_nv525_ | new_nv432_ | new_nv394_;
  assign new_nv440_ = new_n_n198_ & new_n_n67_ & new_nv421_;
  assign new_n_n19_ = new_nv501_ | new_nv553_ | new_nv534_ | new_nv450_ | new_nv403_;
  assign new_nv484_ = new_n_n266_ & new_n_n67_ & new_nv421_;
  assign new_nv496_ = new_n_n241_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv507_ = new_n_n195_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv523_ = new_n_n197_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv534_ = new_n_n232_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv541_ = new_n_n269_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv553_ = new_nv552_ & new_nv421_ & new_nv519_ & new_nv486_;
  assign new_nv578_ = new_n_n34_ & new_nv572_ & new_n_n277_ & new_nv576_;
  assign new_nv604_ = new_n_n39_ & new_nv706_ & new_nv600_;
  assign new_nv612_ = new_n_n38_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_n_n137_ = new_nv654_ | new_nv651_ | new_nv659_ | new_nv656_ | new_nv645_ | new_nv661_ | new_nv648_;
  assign new_nv669_ = new_n_n47_ & new_nv732_ & new_nv699_;
  assign new_nv678_ = new_n_n48_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv693_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n197_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv721_ = new_n_n59_ & new_nv697_;
  assign new_n_n132_ = new_nv767_ | new_nv750_ | new_nv800_ | new_nv783_ | new_nv716_ | new_nv816_ | new_nv733_;
  assign new_nv737_ = new_n_n60_ & new_nv732_ & new_nv699_;
  assign new_n_n123_ = new_nv776_ | new_nv759_ | new_nv809_ | new_nv792_ | new_nv725_ | new_nv825_ | new_nv742_;
  assign new_nv767_ = new_n_n64_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv778_ = new_n_n53_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv786_ = new_n_n277_ & new_n_n61_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv797_ = new_n_n277_ & new_n_n50_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv814_ = new_nv799_ & new_nv627_ & new_n_n157_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv826_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n205_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv834_ = new_n_n31_ & new_nv831_;
  assign new_nv845_ = new_n_n20_ & new_nv831_;
  assign new_n_n114_ = new_nv937_ | new_nv903_ | new_nv1004_ | new_nv971_ | new_nv835_ | new_nv1037_ | new_nv869_;
  assign new_nv875_ = new_n_n24_ & new_nv865_ & new_nv864_;
  assign new_n_n105_ = new_nv946_ | new_nv912_ | new_nv1013_ | new_nv980_ | new_nv844_ | new_nv1046_ | new_nv878_;
  assign new_nv884_ = new_n_n15_ & new_nv865_ & new_nv864_;
  assign new_n_n92_ = new_nv959_ | new_nv925_ | new_nv1026_ | new_nv993_ | new_nv857_ | new_nv1059_ | new_nv891_;
  assign new_nv897_ = new_n_n2_ & new_nv865_ & new_nv864_;
  assign new_nv905_ = new_n_n28_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv916_ = new_n_n17_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv944_ = new_n_n23_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv955_ = new_n_n12_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv975_ = new_nv967_ & new_n_n26_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv990_ = new_nv967_ & new_n_n11_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1002_ = new_n_n277_ & new_nv966_ & new_n_n32_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1009_ = new_n_n277_ & new_nv966_ & new_n_n25_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1020_ = new_n_n277_ & new_nv966_ & new_n_n14_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1047_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n158_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1058_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n184_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1089_ = new_n_n210_ & new_nv1083_ & new_nv1082_;
  assign new_n_n75_ = new_nv1110_ | new_nv1129_ | new_nv1117_ | new_nv1094_ | new_nv1077_;
  assign new_nv1098_ = new_n_n201_ & new_nv1083_ & new_nv1082_;
  assign new_nv1109_ = new_n_n206_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv224_ = new_nv1316_ & new_n_n281_ & new_n_n274_;
  assign new_n_n65_ = new_nv231_ | new_nv230_;
  assign new_nv282_ = new_n_n258_ & new_n_n67_ & new_nv421_;
  assign new_n_n53_ = new_nv335_ | new_nv553_ | new_nv367_ | new_nv290_ | new_nv247_;
  assign new_nv308_ = new_n_n245_ & new_n_n67_ & new_nv421_;
  assign new_n_n39_ = new_nv261_ | new_nv501_ | new_nv553_ | new_nv381_;
  assign new_nv327_ = new_n_n259_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv336_ = new_n_n250_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv394_ = new_n_n210_ & new_n_n68_;
  assign new_nv396_ = new_n_n208_ & new_n_n68_;
  assign new_nv405_ = new_n_n199_ & new_n_n68_;
  assign new_n_n33_ = new_nv487_ | new_nv553_ | new_nv520_ | new_nv422_ | new_nv389_;
  assign new_nv432_ = new_n_n202_ & new_n_n67_ & new_nv421_;
  assign new_n_n24_ = new_nv496_ | new_nv553_ | new_nv529_ | new_nv440_ | new_nv398_;
  assign new_nv450_ = new_n_n239_ & new_n_n67_ & new_nv421_;
  assign new_n_n2_ = new_nv518_ | new_nv553_ | new_nv551_ | new_nv484_ | new_nv420_;
  assign new_nv495_ = new_n_n196_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv497_ = new_n_n240_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv524_ = new_n_n196_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv533_ = new_n_n233_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv542_ = new_n_n268_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv551_ = new_n_n259_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv596_ = new_n_n39_ & new_nv631_;
  assign new_n_n144_ = new_nv596_ | new_nv611_ | new_nv604_ | new_nv618_;
  assign new_nv611_ = new_n_n39_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_nv651_ = new_n_n45_ & new_nv646_ & new_nv749_ & new_nv649_;
  assign new_n_n136_ = new_nv678_ | new_nv673_ | new_nv687_ | new_nv682_ | new_nv663_ | new_nv691_ | new_nv668_;
  assign new_nv679_ = new_n_n47_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv692_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n198_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv722_ = new_n_n58_ & new_nv697_;
  assign new_nv733_ = new_n_n64_ & new_nv732_ & new_nv699_;
  assign new_n_n128_ = new_nv771_ | new_nv754_ | new_nv804_ | new_nv787_ | new_nv720_ | new_nv820_ | new_nv737_;
  assign new_nv742_ = new_n_n55_ & new_nv732_ & new_nv699_;
  assign new_nv768_ = new_n_n63_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv777_ = new_n_n54_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv787_ = new_n_n277_ & new_n_n60_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv796_ = new_n_n277_ & new_n_n51_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv816_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n215_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv825_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n206_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv835_ = new_n_n30_ & new_nv831_;
  assign new_nv844_ = new_n_n21_ & new_nv831_;
  assign new_nv870_ = new_n_n29_ & new_nv865_ & new_nv864_;
  assign new_n_n109_ = new_nv942_ | new_nv908_ | new_nv1009_ | new_nv976_ | new_nv840_ | new_nv1042_ | new_nv874_;
  assign new_nv879_ = new_n_n20_ & new_nv865_ & new_nv864_;
  assign new_n_n100_ = new_nv951_ | new_nv917_ | new_nv1018_ | new_nv985_ | new_nv849_ | new_nv1051_ | new_nv883_;
  assign new_nv892_ = new_n_n7_ & new_nv865_ & new_nv864_;
  assign new_n_n87_ = new_nv964_ | new_nv930_ | new_nv1031_ | new_nv998_ | new_nv862_ | new_nv1064_ | new_nv896_;
  assign new_nv906_ = new_n_n27_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv915_ = new_n_n18_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv945_ = new_n_n22_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv954_ = new_n_n13_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv963_ = new_n_n4_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv991_ = new_nv967_ & new_n_n10_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1001_ = new_n_n277_ & new_nv966_ & new_n_n33_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1010_ = new_n_n277_ & new_nv966_ & new_n_n24_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1019_ = new_n_n277_ & new_nv966_ & new_n_n15_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1048_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n157_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1057_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n185_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_n_n80_ = new_nv1105_ | new_nv1124_ | new_nv1117_ | new_nv1089_ | new_nv1072_;
  assign new_nv1094_ = new_n_n205_ & new_nv1083_ & new_nv1082_;
  assign new_n_n71_ = new_nv1114_ | new_nv1133_ | new_nv1117_ | new_nv1098_ | new_nv1081_;
  assign new_nv1108_ = new_n_n207_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv219_ = new_nv1316_ & new_nv1276_ & new_nv1288_;
  assign new_n_n66_ = new_nv228_ | new_nv226_ | new_nv229_;
  assign new_n_n55_ = new_nv333_ | new_nv553_ | new_nv365_ | new_nv286_ | new_nv245_;
  assign new_nv298_ = new_n_n250_ & new_n_n67_ & new_nv421_;
  assign new_n_n48_ = new_nv340_ | new_nv553_ | new_nv372_ | new_nv300_ | new_nv252_;
  assign new_nv312_ = new_n_n243_ & new_n_n67_ & new_nv421_;
  assign new_nv324_ = new_n_n262_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv335_ = new_n_n251_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv401_ = new_n_n203_ & new_n_n68_;
  assign new_nv412_ = new_n_n238_ & new_n_n68_;
  assign new_nv415_ = new_n_n235_ & new_n_n68_;
  assign new_n_n31_ = new_nv489_ | new_nv553_ | new_nv522_ | new_nv426_ | new_nv391_;
  assign new_nv438_ = new_n_n199_ & new_n_n67_ & new_nv421_;
  assign new_n_n20_ = new_nv500_ | new_nv553_ | new_nv533_ | new_nv448_ | new_nv402_;
  assign new_nv502_ = new_n_n235_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv513_ = new_n_n268_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv528_ = new_n_n238_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv539_ = new_n_n271_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv550_ = new_n_n260_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv619_ = new_nv1316_ & new_n_n182_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_n_n139_ = new_nv632_ | new_nv639_ | new_nv636_ | new_nv642_;
  assign new_nv674_ = new_n_n47_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv691_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n199_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_n_n120_ = new_nv779_ | new_nv762_ | new_nv812_ | new_nv795_ | new_nv728_ | new_nv828_ | new_nv745_;
  assign new_nv756_ = new_n_n58_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv795_ = new_n_n277_ & new_n_n52_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv817_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n214_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv851_ = new_n_n14_ & new_nv831_;
  assign new_nv862_ = new_n_n3_ & new_nv831_;
  assign new_n_n91_ = new_nv960_ | new_nv926_ | new_nv1027_ | new_nv994_ | new_nv858_ | new_nv1060_ | new_nv892_;
  assign new_nv900_ = new_n_n33_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv922_ = new_n_n11_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv935_ = new_n_n32_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv992_ = new_nv967_ & new_n_n9_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1004_ = new_n_n277_ & new_nv966_ & new_n_n30_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1015_ = new_n_n277_ & new_nv966_ & new_n_n19_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1026_ = new_n_n277_ & new_nv966_ & new_n_n8_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1038_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n167_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1090_ = new_n_n209_ & new_nv1083_ & new_nv1082_;
  assign new_n_n74_ = new_nv1111_ | new_nv1130_ | new_nv1117_ | new_nv1095_ | new_nv1078_;
  assign new_nv1104_ = new_n_n211_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv1117_ = new_nv1116_ & new_nv1082_ & new_nv1316_ & new_nv1099_;
  assign new_nv582_ = ~new_nv1143_;
  assign new_nv222_ = new_nv1316_ & new_n_n281_ & new_nv1288_ & new_nv1295_ & new_nv1289_;
  assign new_n_n67_ = new_nv224_ | new_nv219_ | new_nv222_ | new_nv223_;
  assign new_nv288_ = new_n_n255_ & new_n_n67_ & new_nv421_;
  assign new_n_n50_ = new_nv338_ | new_nv553_ | new_nv370_ | new_nv296_ | new_nv250_;
  assign new_nv302_ = new_n_n248_ & new_n_n67_ & new_nv421_;
  assign new_n_n43_ = new_nv497_ | new_nv553_ | new_nv377_ | new_nv310_ | new_nv257_;
  assign new_nv325_ = new_n_n261_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv334_ = new_n_n252_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv402_ = new_n_n202_ & new_n_n68_;
  assign new_nv411_ = new_n_n239_ & new_n_n68_;
  assign new_nv416_ = new_n_n234_ & new_n_n68_;
  assign new_nv426_ = new_n_n205_ & new_n_n67_ & new_nv421_;
  assign new_n_n25_ = new_nv495_ | new_nv553_ | new_nv528_ | new_nv438_ | new_nv397_;
  assign new_nv448_ = new_n_n240_ & new_n_n67_ & new_nv421_;
  assign new_nv503_ = new_n_n234_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv512_ = new_n_n269_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv517_ = new_n_n264_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv540_ = new_n_n270_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv549_ = new_n_n261_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv620_ = new_nv1316_ & new_n_n181_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_nv636_ = new_n_n44_ & new_nv706_ & new_nv600_;
  assign new_nv675_ = new_n_n46_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv689_ = new_nv799_ & new_nv627_ & new_n_n173_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv746_ = new_n_n51_ & new_nv732_ & new_nv699_;
  assign new_nv755_ = new_n_n59_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv785_ = new_n_n277_ & new_n_n62_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv827_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n204_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv852_ = new_n_n13_ & new_nv831_;
  assign new_nv861_ = new_n_n4_ & new_nv831_;
  assign new_nv893_ = new_n_n6_ & new_nv865_ & new_nv864_;
  assign new_n_n86_ = new_nv965_ | new_nv931_ | new_nv1032_ | new_nv999_ | new_nv863_ | new_nv1065_ | new_nv897_;
  assign new_nv923_ = new_n_n10_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv934_ = new_n_n33_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv993_ = new_nv967_ & new_n_n8_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1003_ = new_n_n277_ & new_nv966_ & new_n_n31_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1025_ = new_n_n277_ & new_nv966_ & new_n_n9_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1027_ = new_n_n277_ & new_nv966_ & new_n_n7_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1037_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n168_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_n_n79_ = new_nv1106_ | new_nv1125_ | new_nv1117_ | new_nv1090_ | new_nv1073_;
  assign new_nv1095_ = new_n_n204_ & new_nv1083_ & new_nv1082_;
  assign new_nv1105_ = new_n_n210_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv1114_ = new_n_n201_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_n_n68_ = new_n_n277_ | new_nv215_;
  assign new_n_n56_ = new_nv332_ | new_nv553_ | new_nv364_ | new_nv284_ | new_nv244_;
  assign new_nv296_ = new_n_n251_ & new_n_n67_ & new_nv421_;
  assign new_n_n47_ = new_nv341_ | new_nv553_ | new_nv373_ | new_nv302_ | new_nv253_;
  assign new_nv314_ = new_n_n242_ & new_n_n67_ & new_nv421_;
  assign new_n_n35_ = new_nv265_ | new_nv505_ | new_nv553_ | new_nv385_;
  assign new_nv333_ = new_n_n253_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv399_ = new_n_n205_ & new_n_n68_;
  assign new_nv410_ = new_n_n240_ & new_n_n68_;
  assign new_nv417_ = new_n_n233_ & new_n_n68_;
  assign new_n_n30_ = new_nv490_ | new_nv553_ | new_nv523_ | new_nv428_ | new_nv392_;
  assign new_nv436_ = new_n_n200_ & new_n_n67_ & new_nv421_;
  assign new_n_n21_ = new_nv499_ | new_nv553_ | new_nv532_ | new_nv446_ | new_nv401_;
  assign new_nv500_ = new_n_n237_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv511_ = new_n_n270_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv518_ = new_n_n263_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv530_ = new_n_n236_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv548_ = new_n_n262_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv617_ = new_nv1316_ & new_n_n184_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_nv633_ = new_n_n43_ & new_nv631_;
  assign new_nv642_ = new_nv1316_ & new_n_n178_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_nv664_ = new_n_n47_ & new_nv697_;
  assign new_n_n121_ = new_nv778_ | new_nv761_ | new_nv811_ | new_nv794_ | new_nv727_ | new_nv827_ | new_nv744_;
  assign new_nv754_ = new_n_n60_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv774_ = new_n_n57_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv838_ = new_n_n27_ & new_nv831_;
  assign new_nv849_ = new_n_n16_ & new_nv831_;
  assign new_nv860_ = new_n_n5_ & new_nv831_;
  assign new_nv909_ = new_n_n24_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv920_ = new_n_n13_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv931_ = new_n_n2_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv994_ = new_nv967_ & new_n_n7_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1013_ = new_n_n277_ & new_nv966_ & new_n_n21_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1024_ = new_n_n277_ & new_nv966_ & new_n_n10_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1091_ = new_n_n208_ & new_nv1083_ & new_nv1082_;
  assign new_n_n73_ = new_nv1112_ | new_nv1131_ | new_nv1117_ | new_nv1096_ | new_nv1079_;
  assign new_nv1102_ = new_n_n213_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv1113_ = new_n_n202_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv215_ = new_n_n282_ & new_n_n281_ & new_n_n280_;
  assign new_nv231_ = new_nv1316_ & new_nv1309_ & new_n_n275_ & new_nv1295_;
  assign new_nv286_ = new_n_n256_ & new_n_n67_ & new_nv421_;
  assign new_n_n51_ = new_nv337_ | new_nv553_ | new_nv369_ | new_nv294_ | new_nv249_;
  assign new_nv304_ = new_n_n247_ & new_n_n67_ & new_nv421_;
  assign new_n_n42_ = new_nv498_ | new_nv553_ | new_nv378_ | new_nv312_ | new_nv258_;
  assign new_n_n34_ = new_nv266_ | new_nv506_ | new_nv553_ | new_nv386_;
  assign new_nv332_ = new_n_n254_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv400_ = new_n_n204_ & new_n_n68_;
  assign new_nv409_ = new_n_n241_ & new_n_n68_;
  assign new_nv418_ = new_n_n232_ & new_n_n68_;
  assign new_nv428_ = new_n_n204_ & new_n_n67_ & new_nv421_;
  assign new_n_n26_ = new_nv494_ | new_nv553_ | new_nv527_ | new_nv436_ | new_nv396_;
  assign new_nv446_ = new_n_n241_ & new_n_n67_ & new_nv421_;
  assign new_nv501_ = new_n_n236_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv510_ = new_n_n271_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv520_ = new_n_n200_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv529_ = new_n_n237_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv538_ = new_n_n272_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv618_ = new_nv1316_ & new_n_n183_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_nv632_ = new_n_n44_ & new_nv631_;
  assign new_nv643_ = new_nv1316_ & new_n_n177_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_nv663_ = new_n_n48_ & new_nv697_;
  assign new_nv745_ = new_n_n52_ & new_nv732_ & new_nv699_;
  assign new_nv753_ = new_n_n61_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv762_ = new_n_n52_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv848_ = new_n_n17_ & new_nv831_;
  assign new_nv850_ = new_n_n15_ & new_nv831_;
  assign new_nv859_ = new_n_n6_ & new_nv831_;
  assign new_nv910_ = new_n_n23_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv919_ = new_n_n14_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv921_ = new_n_n12_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv1005_ = new_n_n277_ & new_nv966_ & new_n_n29_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1014_ = new_n_n277_ & new_nv966_ & new_n_n20_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1023_ = new_n_n277_ & new_nv966_ & new_n_n11_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_n_n78_ = new_nv1107_ | new_nv1126_ | new_nv1117_ | new_nv1091_ | new_nv1074_;
  assign new_nv1096_ = new_n_n203_ & new_nv1083_ & new_nv1082_;
  assign new_nv1103_ = new_n_n212_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv1112_ = new_n_n203_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv241_ = new_n_n268_ & new_n_n68_;
  assign new_nv252_ = new_n_n257_ & new_n_n68_;
  assign new_nv263_ = new_n_n246_ & new_n_n68_;
  assign new_n_n61_ = new_nv327_ | new_nv553_ | new_nv359_ | new_nv274_ | new_nv239_;
  assign new_nv342_ = new_n_n244_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv365_ = new_n_n249_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv376_ = new_n_n226_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv389_ = new_n_n215_ & new_n_n68_;
  assign new_nv456_ = new_n_n236_ & new_n_n67_ & new_nv421_;
  assign new_n_n11_ = new_nv509_ | new_nv553_ | new_nv542_ | new_nv466_ | new_nv411_;
  assign new_nv478_ = new_n_n269_ & new_n_n67_ & new_nv421_;
  assign new_nv490_ = new_n_n201_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv506_ = new_n_n231_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv581_ = new_n_n191_ & new_nv572_ & new_nv1316_ & new_nv576_ & new_nv1143_;
  assign new_nv598_ = new_n_n37_ & new_nv631_;
  assign new_n_n142_ = new_nv598_ | new_nv613_ | new_nv606_ | new_nv620_;
  assign new_nv626_ = new_n_n42_ & new_nv706_ & new_nv624_;
  assign new_nv640_ = new_n_n43_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_nv734_ = new_n_n63_ & new_nv732_ & new_nv699_;
  assign new_n_n126_ = new_nv773_ | new_nv756_ | new_nv806_ | new_nv789_ | new_nv722_ | new_nv822_ | new_nv739_;
  assign new_n_n118_ = new_nv781_ | new_nv764_ | new_nv814_ | new_nv797_ | new_nv730_ | new_nv830_ | new_nv747_;
  assign new_nv760_ = new_n_n54_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv773_ = new_n_n58_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv839_ = new_n_n26_ & new_nv831_;
  assign new_nv855_ = new_n_n10_ & new_nv831_;
  assign new_nv867_ = new_n_n32_ & new_nv865_ & new_nv864_;
  assign new_n_n111_ = new_nv940_ | new_nv906_ | new_nv1007_ | new_nv974_ | new_nv838_ | new_nv1040_ | new_nv872_;
  assign new_nv878_ = new_n_n21_ & new_nv865_ & new_nv864_;
  assign new_nv926_ = new_n_n7_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv939_ = new_n_n28_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv950_ = new_n_n17_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv961_ = new_n_n6_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv974_ = new_nv967_ & new_n_n27_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1030_ = new_n_n277_ & new_nv966_ & new_n_n4_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1042_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n163_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1053_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n176_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1064_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n186_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1076_ = new_n_n206_ & new_nv1066_;
  assign new_n_n83_ = new_nv1102_ | new_nv1121_ | new_nv1117_ | new_nv1086_ | new_nv1069_;
  assign new_nv559_ = ~new_nv557_;
  assign new_nv242_ = new_n_n267_ & new_n_n68_;
  assign new_nv251_ = new_n_n258_ & new_n_n68_;
  assign new_nv264_ = new_n_n245_ & new_n_n68_;
  assign new_nv274_ = new_n_n262_ & new_n_n67_ & new_nv421_;
  assign new_nv343_ = new_n_n243_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv364_ = new_n_n250_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv377_ = new_n_n225_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv386_ = new_n_n216_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_n_n16_ = new_nv504_ | new_nv553_ | new_nv537_ | new_nv456_ | new_nv406_;
  assign new_nv466_ = new_n_n231_ & new_n_n67_ & new_nv421_;
  assign new_n_n5_ = new_nv515_ | new_nv553_ | new_nv548_ | new_nv478_ | new_nv417_;
  assign new_nv489_ = new_n_n202_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv516_ = new_n_n265_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv566_ = new_n_n277_ & new_n_n195_ & new_nv559_ & new_nv660_ & new_nv556_ & new_nv562_;
  assign new_nv599_ = new_n_n36_ & new_nv631_;
  assign new_nv606_ = new_n_n37_ & new_nv706_ & new_nv600_;
  assign new_n_n140_ = new_nv623_ | new_nv628_ | new_nv626_ | new_nv630_;
  assign new_nv639_ = new_n_n44_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_n_n131_ = new_nv768_ | new_nv751_ | new_nv801_ | new_nv784_ | new_nv717_ | new_nv817_ | new_nv734_;
  assign new_nv739_ = new_n_n58_ & new_nv732_ & new_nv699_;
  assign new_nv750_ = new_n_n64_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv759_ = new_n_n55_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv784_ = new_n_n277_ & new_n_n63_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv828_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n203_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv856_ = new_n_n9_ & new_nv831_;
  assign new_n_n117_ = new_nv934_ | new_nv900_ | new_nv1001_ | new_nv968_ | new_nv832_ | new_nv1034_ | new_nv866_;
  assign new_nv873_ = new_n_n26_ & new_nv865_ & new_nv864_;
  assign new_n_n106_ = new_nv945_ | new_nv911_ | new_nv1012_ | new_nv979_ | new_nv843_ | new_nv1045_ | new_nv877_;
  assign new_nv927_ = new_n_n6_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv938_ = new_n_n29_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv951_ = new_n_n16_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv960_ = new_n_n7_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv984_ = new_nv967_ & new_n_n17_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1031_ = new_n_n277_ & new_nv966_ & new_n_n3_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1041_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n164_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1054_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n178_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1063_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n188_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1077_ = new_n_n205_ & new_nv1066_;
  assign new_nv1086_ = new_n_n213_ & new_nv1083_ & new_nv1082_;
  assign new_nv562_ = ~new_nv560_;
  assign new_nv243_ = new_n_n266_ & new_n_n68_;
  assign new_nv254_ = new_n_n255_ & new_n_n68_;
  assign new_nv261_ = new_n_n248_ & new_n_n68_;
  assign new_n_n62_ = new_nv326_ | new_nv553_ | new_nv358_ | new_nv272_ | new_nv238_;
  assign new_n_n54_ = new_nv334_ | new_nv553_ | new_nv366_ | new_nv288_ | new_nv246_;
  assign new_nv356_ = new_n_n258_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv367_ = new_n_n247_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv374_ = new_n_n228_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv385_ = new_n_n217_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv403_ = new_n_n201_ & new_n_n68_;
  assign new_nv414_ = new_n_n236_ & new_n_n68_;
  assign new_nv458_ = new_n_n235_ & new_n_n67_ & new_nv421_;
  assign new_n_n10_ = new_nv510_ | new_nv553_ | new_nv543_ | new_nv468_ | new_nv412_;
  assign new_nv476_ = new_n_n270_ & new_n_n67_ & new_nv421_;
  assign new_nv488_ = new_n_n203_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv504_ = new_n_n233_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv515_ = new_n_n266_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv568_ = new_nv1316_ & new_nv556_ & new_nv562_ & new_nv559_ & new_nv660_;
  assign new_nv585_ = new_nv1146_ & new_n_n189_ & new_nv576_ & new_nv582_ & new_nv572_ & new_nv1316_;
  assign new_n_n143_ = new_nv597_ | new_nv612_ | new_nv605_ | new_nv619_;
  assign new_nv621_ = new_nv1316_ & new_n_n180_ & new_nv600_ & new_nv1316_ & new_nv627_ & new_n_n187_;
  assign new_n_n138_ = new_nv633_ | new_nv640_ | new_nv637_ | new_nv643_;
  assign new_nv709_ = new_n_n277_ & new_nv652_ & new_n_n49_ & new_nv649_ & new_nv627_ & new_nv696_ & new_nv699_;
  assign new_nv724_ = new_n_n56_ & new_nv697_;
  assign new_n_n119_ = new_nv780_ | new_nv763_ | new_nv813_ | new_nv796_ | new_nv729_ | new_nv829_ | new_nv746_;
  assign new_nv758_ = new_n_n56_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv794_ = new_n_n277_ & new_n_n53_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv818_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n213_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv853_ = new_n_n12_ & new_nv831_;
  assign new_nv866_ = new_n_n33_ & new_nv865_ & new_nv864_;
  assign new_n_n101_ = new_nv950_ | new_nv916_ | new_nv1017_ | new_nv984_ | new_nv848_ | new_nv1050_ | new_nv882_;
  assign new_nv888_ = new_n_n11_ & new_nv865_ & new_nv864_;
  assign new_nv924_ = new_n_n9_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv937_ = new_n_n30_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv952_ = new_n_n15_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv972_ = new_nv967_ & new_n_n29_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv983_ = new_nv967_ & new_n_n18_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1028_ = new_n_n277_ & new_nv966_ & new_n_n6_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1040_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n165_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1055_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n177_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1067_ = new_n_n215_ & new_nv1066_;
  assign new_nv1074_ = new_n_n208_ & new_nv1066_;
  assign new_n_n84_ = new_nv1101_ | new_nv1120_ | new_nv1117_ | new_nv1085_ | new_nv1068_;
  assign new_nv572_ = ~new_nv569_;
  assign new_nv244_ = new_n_n265_ & new_n_n68_;
  assign new_nv253_ = new_n_n256_ & new_n_n68_;
  assign new_nv262_ = new_n_n247_ & new_n_n68_;
  assign new_nv272_ = new_n_n263_ & new_n_n67_ & new_nv421_;
  assign new_n_n49_ = new_nv339_ | new_nv553_ | new_nv371_ | new_nv298_ | new_nv251_;
  assign new_nv357_ = new_n_n257_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv366_ = new_n_n248_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv375_ = new_n_n227_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv384_ = new_n_n218_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv404_ = new_n_n200_ & new_n_n68_;
  assign new_nv413_ = new_n_n237_ & new_n_n68_;
  assign new_n_n15_ = new_nv505_ | new_nv553_ | new_nv538_ | new_nv458_ | new_nv407_;
  assign new_nv468_ = new_n_n195_ & new_n_n67_ & new_nv421_;
  assign new_n_n6_ = new_nv514_ | new_nv553_ | new_nv547_ | new_nv476_ | new_nv416_;
  assign new_nv487_ = new_n_n204_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv505_ = new_n_n232_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv514_ = new_n_n267_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv570_ = new_n_n35_ & new_nv569_;
  assign new_nv584_ = new_nv1146_ & new_n_n190_ & new_nv576_ & new_nv582_ & new_nv572_ & new_nv1316_;
  assign new_nv597_ = new_n_n38_ & new_nv631_;
  assign new_nv623_ = new_n_n42_ & new_nv622_;
  assign new_nv637_ = new_n_n43_ & new_nv706_ & new_nv600_;
  assign new_nv712_ = new_nv627_ & new_nv649_ & new_nv799_ & new_n_n172_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv696_;
  assign new_nv723_ = new_n_n57_ & new_nv697_;
  assign new_nv747_ = new_n_n50_ & new_nv732_ & new_nv699_;
  assign new_nv757_ = new_n_n57_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv806_ = new_nv799_ & new_nv627_ & new_n_n165_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv807_ = new_nv799_ & new_nv627_ & new_n_n164_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv854_ = new_n_n11_ & new_nv831_;
  assign new_nv863_ = new_n_n2_ & new_nv831_;
  assign new_nv883_ = new_n_n16_ & new_nv865_ & new_nv864_;
  assign new_n_n96_ = new_nv955_ | new_nv921_ | new_nv1022_ | new_nv989_ | new_nv853_ | new_nv1055_ | new_nv887_;
  assign new_nv925_ = new_n_n8_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv936_ = new_n_n31_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv962_ = new_n_n5_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv973_ = new_nv967_ & new_n_n28_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv982_ = new_nv967_ & new_n_n19_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1029_ = new_n_n277_ & new_nv966_ & new_n_n5_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1039_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n166_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1056_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n179_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1065_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n192_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1075_ = new_n_n207_ & new_nv1066_;
  assign new_nv1085_ = new_n_n214_ & new_nv1083_ & new_nv1082_;
  assign new_nv576_ = ~new_nv573_;
  assign new_nv245_ = new_n_n264_ & new_n_n68_;
  assign new_nv256_ = new_n_n253_ & new_n_n68_;
  assign new_nv268_ = new_n_n265_ & new_n_n67_ & new_nv421_;
  assign new_n_n59_ = new_nv329_ | new_nv553_ | new_nv361_ | new_nv278_ | new_nv241_;
  assign new_n_n44_ = new_nv496_ | new_nv553_ | new_nv376_ | new_nv308_ | new_nv256_;
  assign new_nv358_ = new_n_n256_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv369_ = new_n_n245_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv380_ = new_n_n222_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv393_ = new_n_n211_ & new_n_n68_;
  assign new_nv424_ = new_n_n206_ & new_n_n67_ & new_nv421_;
  assign new_n_n27_ = new_nv493_ | new_nv553_ | new_nv526_ | new_nv434_ | new_nv395_;
  assign new_nv460_ = new_n_n234_ & new_n_n67_ & new_nv421_;
  assign new_n_n9_ = new_nv511_ | new_nv553_ | new_nv544_ | new_nv470_ | new_nv413_;
  assign new_nv482_ = new_n_n267_ & new_n_n67_ & new_nv421_;
  assign new_nv494_ = new_n_n197_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv525_ = new_n_n241_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv536_ = new_n_n195_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv547_ = new_n_n263_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv571_ = new_n_n34_ & new_nv569_;
  assign new_nv589_ = new_nv587_ & new_nv582_ & new_n_n189_ & new_nv1316_ & new_nv586_ & new_nv572_ & new_nv576_;
  assign new_nv603_ = new_n_n40_ & new_nv706_ & new_nv600_;
  assign new_nv610_ = new_n_n40_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_nv654_ = new_n_n45_ & new_nv646_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv670_ = new_n_n46_ & new_nv732_ & new_nv699_;
  assign new_nv687_ = new_nv799_ & new_nv627_ & new_n_n175_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv707_ = new_nv706_ & new_n_n49_ & new_nv699_ & new_nv652_ & new_nv696_ & new_nv649_;
  assign new_nv714_ = new_nv652_ & new_nv699_ & new_nv1310_ & new_nv1316_ & new_nv1315_ & new_nv1263_ & new_nv1287_ & new_nv1316_ & new_n_n281_ & new_n_n280_ & new_n_n200_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv696_;
  assign new_nv726_ = new_n_n54_ & new_nv697_;
  assign new_nv736_ = new_n_n61_ & new_nv732_ & new_nv699_;
  assign new_n_n124_ = new_nv775_ | new_nv758_ | new_nv808_ | new_nv791_ | new_nv724_ | new_nv824_ | new_nv741_;
  assign new_nv769_ = new_n_n62_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv780_ = new_n_n51_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv792_ = new_n_n277_ & new_n_n55_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv805_ = new_nv799_ & new_nv627_ & new_n_n166_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv808_ = new_nv799_ & new_nv627_ & new_n_n163_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv820_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n211_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv832_ = new_n_n33_ & new_nv831_;
  assign new_nv843_ = new_n_n22_ & new_nv831_;
  assign new_n_n113_ = new_nv938_ | new_nv904_ | new_nv1005_ | new_nv972_ | new_nv836_ | new_nv1038_ | new_nv870_;
  assign new_nv876_ = new_n_n23_ & new_nv865_ & new_nv864_;
  assign new_n_n102_ = new_nv949_ | new_nv915_ | new_nv1016_ | new_nv983_ | new_nv847_ | new_nv1049_ | new_nv881_;
  assign new_nv887_ = new_n_n12_ & new_nv865_ & new_nv864_;
  assign new_n_n95_ = new_nv956_ | new_nv922_ | new_nv1023_ | new_nv990_ | new_nv854_ | new_nv1056_ | new_nv888_;
  assign new_nv894_ = new_n_n5_ & new_nv865_ & new_nv864_;
  assign new_nv903_ = new_n_n30_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv914_ = new_n_n19_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv930_ = new_n_n3_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv946_ = new_n_n21_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv957_ = new_n_n10_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv970_ = new_nv967_ & new_n_n31_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv981_ = new_nv967_ & new_n_n20_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv995_ = new_nv967_ & new_n_n6_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1007_ = new_n_n277_ & new_nv966_ & new_n_n27_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1018_ = new_n_n277_ & new_nv966_ & new_n_n16_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1035_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n170_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1046_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n159_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1049_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n172_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1060_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n182_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1072_ = new_n_n210_ & new_nv1066_;
  assign new_n_n85_ = new_nv1100_ | new_nv1119_ | new_nv1117_ | new_nv1084_ | new_nv1067_;
  assign new_nv1097_ = new_n_n202_ & new_nv1083_ & new_nv1082_;
  assign new_nv1107_ = new_n_n208_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv486_ = ~new_n_n67_;
  assign new_nv246_ = new_n_n263_ & new_n_n68_;
  assign new_nv255_ = new_n_n254_ & new_n_n68_;
  assign new_n_n64_ = new_nv324_ | new_nv553_ | new_nv356_ | new_nv268_ | new_nv236_;
  assign new_nv278_ = new_n_n260_ & new_n_n67_ & new_nv421_;
  assign new_n_n37_ = new_nv263_ | new_nv503_ | new_nv553_ | new_nv383_;
  assign new_nv359_ = new_n_n255_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv368_ = new_n_n246_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv381_ = new_n_n221_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv392_ = new_n_n212_ & new_n_n68_;
  assign new_n_n32_ = new_nv488_ | new_nv553_ | new_nv521_ | new_nv424_ | new_nv390_;
  assign new_nv434_ = new_n_n201_ & new_n_n67_ & new_nv421_;
  assign new_n_n14_ = new_nv506_ | new_nv553_ | new_nv539_ | new_nv460_ | new_nv408_;
  assign new_nv470_ = new_n_n273_ & new_n_n67_ & new_nv421_;
  assign new_n_n3_ = new_nv517_ | new_nv553_ | new_nv550_ | new_nv482_ | new_nv419_;
  assign new_nv493_ = new_n_n198_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv526_ = new_n_n240_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv535_ = new_n_n231_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv564_ = new_n_n192_ & new_nv556_ & new_nv562_ & new_nv559_ & new_nv799_;
  assign new_nv574_ = new_n_n35_ & new_nv573_ & new_nv572_;
  assign new_nv588_ = new_nv587_ & new_nv582_ & new_n_n190_ & new_nv1316_ & new_nv586_ & new_nv572_ & new_nv576_;
  assign new_n_n145_ = new_nv595_ | new_nv610_ | new_nv603_ | new_nv617_;
  assign new_nv609_ = new_n_n41_ & new_nv600_ & new_n_n277_ & new_nv627_;
  assign new_nv656_ = new_n_n277_ & new_n_n45_ & new_nv649_ & new_nv627_ & new_nv646_ & new_nv652_;
  assign new_n_n135_ = new_nv679_ | new_nv674_ | new_nv688_ | new_nv683_ | new_nv664_ | new_nv692_ | new_nv669_;
  assign new_nv688_ = new_nv799_ & new_nv627_ & new_n_n174_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv704_ = new_n_n49_ & new_nv696_ & new_nv649_ & new_nv699_ & new_nv749_;
  assign new_nv716_ = new_n_n64_ & new_nv697_;
  assign new_nv725_ = new_n_n55_ & new_nv697_;
  assign new_n_n129_ = new_nv770_ | new_nv753_ | new_nv803_ | new_nv786_ | new_nv719_ | new_nv819_ | new_nv736_;
  assign new_nv741_ = new_n_n56_ & new_nv732_ & new_nv699_;
  assign new_nv770_ = new_n_n61_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv779_ = new_n_n52_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv793_ = new_n_n277_ & new_n_n54_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv804_ = new_nv799_ & new_nv627_ & new_n_n167_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv809_ = new_nv799_ & new_nv627_ & new_n_n162_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv819_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n212_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv833_ = new_n_n32_ & new_nv831_;
  assign new_nv842_ = new_n_n23_ & new_nv831_;
  assign new_nv871_ = new_n_n28_ & new_nv865_ & new_nv864_;
  assign new_n_n108_ = new_nv943_ | new_nv909_ | new_nv1010_ | new_nv977_ | new_nv841_ | new_nv1043_ | new_nv875_;
  assign new_nv882_ = new_n_n17_ & new_nv865_ & new_nv864_;
  assign new_n_n97_ = new_nv954_ | new_nv920_ | new_nv1021_ | new_nv988_ | new_nv852_ | new_nv1054_ | new_nv886_;
  assign new_nv889_ = new_n_n10_ & new_nv865_ & new_nv864_;
  assign new_n_n90_ = new_nv961_ | new_nv927_ | new_nv1028_ | new_nv995_ | new_nv859_ | new_nv1061_ | new_nv893_;
  assign new_nv904_ = new_n_n29_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv913_ = new_n_n20_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv942_ = new_n_n25_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv947_ = new_n_n20_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv956_ = new_n_n11_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv971_ = new_nv967_ & new_n_n30_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv980_ = new_nv967_ & new_n_n21_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv985_ = new_nv967_ & new_n_n16_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1008_ = new_n_n277_ & new_nv966_ & new_n_n26_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1017_ = new_n_n277_ & new_nv966_ & new_n_n17_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1036_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n169_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1045_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n160_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1050_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n175_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1059_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n183_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1073_ = new_n_n209_ & new_nv1066_;
  assign new_nv1084_ = new_n_n215_ & new_nv1083_ & new_nv1082_;
  assign new_n_n72_ = new_nv1113_ | new_nv1132_ | new_nv1117_ | new_nv1097_ | new_nv1080_;
  assign new_nv1106_ = new_n_n209_ & new_nv1082_ & new_n_n277_ & new_nv1099_;
  assign new_nv519_ = ~new_n_n66_;
  assign new_nv247_ = new_n_n262_ & new_n_n68_;
  assign new_nv258_ = new_n_n251_ & new_n_n68_;
  assign new_nv265_ = new_n_n244_ & new_n_n68_;
  assign new_n_n60_ = new_nv328_ | new_nv553_ | new_nv360_ | new_nv276_ | new_nv240_;
  assign new_nv330_ = new_n_n256_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv360_ = new_n_n254_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv371_ = new_n_n243_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv378_ = new_n_n224_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv391_ = new_n_n213_ & new_n_n68_;
  assign new_nv444_ = new_n_n196_ & new_n_n67_ & new_nv421_;
  assign new_n_n17_ = new_nv503_ | new_nv553_ | new_nv536_ | new_nv454_ | new_nv405_;
  assign new_nv462_ = new_n_n233_ & new_n_n67_ & new_nv421_;
  assign new_n_n8_ = new_nv512_ | new_nv553_ | new_nv545_ | new_nv472_ | new_nv414_;
  assign new_nv480_ = new_n_n268_ & new_n_n67_ & new_nv421_;
  assign new_nv492_ = new_n_n199_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv527_ = new_n_n239_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv545_ = new_n_n265_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv561_ = new_n_n193_ & new_nv556_ & new_nv560_ & new_nv559_;
  assign new_n_n148_ = new_nv584_ | new_nv577_ | new_nv574_ | new_nv570_ | new_nv591_ | new_nv588_;
  assign new_nv592_ = new_nv586_ & new_nv1316_ & new_nv1316_ & new_n_n187_ & new_n_n186_ & new_nv582_ & new_nv590_ & new_nv576_ & new_nv572_;
  assign new_nv602_ = new_n_n41_ & new_nv706_ & new_nv600_;
  assign new_n_n141_ = new_nv599_ | new_nv614_ | new_nv607_ | new_nv621_;
  assign new_nv659_ = new_nv799_ & new_nv627_ & new_n_n176_ & new_nv652_ & new_nv1316_ & new_nv646_ & new_nv649_;
  assign new_nv673_ = new_n_n48_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv683_ = new_n_n277_ & new_n_n47_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv701_ = new_n_n49_ & new_nv696_ & new_nv732_ & new_nv699_;
  assign new_nv717_ = new_n_n63_ & new_nv697_;
  assign new_nv728_ = new_n_n52_ & new_nv697_;
  assign new_nv735_ = new_n_n62_ & new_nv732_ & new_nv699_;
  assign new_n_n125_ = new_nv774_ | new_nv757_ | new_nv807_ | new_nv790_ | new_nv723_ | new_nv823_ | new_nv740_;
  assign new_nv751_ = new_n_n63_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv771_ = new_n_n60_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv783_ = new_n_n277_ & new_n_n64_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv790_ = new_n_n277_ & new_n_n57_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv803_ = new_nv799_ & new_nv627_ & new_n_n168_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv810_ = new_nv799_ & new_nv627_ & new_n_n161_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv822_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n209_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv829_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n202_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv841_ = new_n_n24_ & new_nv831_;
  assign new_nv857_ = new_n_n8_ & new_nv831_;
  assign new_nv868_ = new_n_n31_ & new_nv865_ & new_nv864_;
  assign new_n_n112_ = new_nv939_ | new_nv905_ | new_nv1006_ | new_nv973_ | new_nv837_ | new_nv1039_ | new_nv871_;
  assign new_nv877_ = new_n_n22_ & new_nv865_ & new_nv864_;
  assign new_n_n103_ = new_nv948_ | new_nv914_ | new_nv1015_ | new_nv982_ | new_nv846_ | new_nv1048_ | new_nv880_;
  assign new_nv886_ = new_n_n13_ & new_nv865_ & new_nv864_;
  assign new_n_n94_ = new_nv957_ | new_nv923_ | new_nv1024_ | new_nv991_ | new_nv855_ | new_nv1057_ | new_nv889_;
  assign new_nv895_ = new_n_n4_ & new_nv865_ & new_nv864_;
  assign new_nv901_ = new_n_n32_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv912_ = new_n_n21_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv928_ = new_n_n5_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv941_ = new_n_n26_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv948_ = new_n_n19_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv959_ = new_n_n8_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv968_ = new_nv967_ & new_n_n33_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv979_ = new_nv967_ & new_n_n22_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv986_ = new_nv967_ & new_n_n15_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv997_ = new_nv967_ & new_n_n4_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1016_ = new_n_n277_ & new_nv966_ & new_n_n18_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1032_ = new_n_n277_ & new_nv966_ & new_n_n2_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1044_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n161_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1051_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n174_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1062_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n180_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1070_ = new_n_n212_ & new_nv1066_;
  assign new_nv1081_ = new_n_n201_ & new_nv1066_;
  assign new_nv1087_ = new_n_n212_ & new_nv1083_ & new_nv1082_;
  assign new_n_n77_ = new_nv1108_ | new_nv1127_ | new_nv1117_ | new_nv1092_ | new_nv1075_;
  assign new_nv552_ = ~new_n_n65_;
  assign new_nv248_ = new_n_n261_ & new_n_n68_;
  assign new_nv257_ = new_n_n252_ & new_n_n68_;
  assign new_nv266_ = new_n_n243_ & new_n_n68_;
  assign new_nv276_ = new_n_n261_ & new_n_n67_ & new_nv421_;
  assign new_nv340_ = new_n_n246_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv361_ = new_n_n253_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv370_ = new_n_n244_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv379_ = new_n_n223_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv390_ = new_n_n214_ & new_n_n68_;
  assign new_n_n22_ = new_nv498_ | new_nv553_ | new_nv531_ | new_nv444_ | new_nv400_;
  assign new_nv454_ = new_n_n237_ & new_n_n67_ & new_nv421_;
  assign new_n_n13_ = new_nv507_ | new_nv553_ | new_nv540_ | new_nv462_ | new_nv409_;
  assign new_nv472_ = new_n_n272_ & new_n_n67_ & new_nv421_;
  assign new_n_n4_ = new_nv516_ | new_nv553_ | new_nv549_ | new_nv480_ | new_nv418_;
  assign new_nv491_ = new_n_n200_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv537_ = new_n_n273_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv546_ = new_n_n264_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_n_n149_ = new_nv566_ | new_nv561_ | new_nv558_ | new_nv555_ | new_nv564_ | new_nv568_;
  assign new_nv575_ = new_n_n34_ & new_nv573_ & new_nv572_;
  assign new_nv591_ = new_nv586_ & new_nv1316_ & new_nv1316_ & new_n_n187_ & new_n_n188_ & new_nv582_ & new_nv590_ & new_nv576_ & new_nv572_;
  assign new_n_n146_ = new_nv594_ | new_nv609_ | new_nv602_ | new_nv616_;
  assign new_nv607_ = new_n_n36_ & new_nv706_ & new_nv600_;
  assign new_nv661_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n196_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv646_;
  assign new_n_n134_ = new_nv680_ | new_nv675_ | new_nv689_ | new_nv684_ | new_nv665_ | new_nv693_ | new_nv670_;
  assign new_nv684_ = new_n_n277_ & new_n_n46_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_n_n133_ = new_nv707_ | new_nv704_ | new_nv712_ | new_nv709_ | new_nv714_ | new_nv695_ | new_nv701_ | new_nv698_;
  assign new_nv718_ = new_n_n62_ & new_nv697_;
  assign new_nv727_ = new_n_n53_ & new_nv697_;
  assign new_n_n130_ = new_nv769_ | new_nv752_ | new_nv802_ | new_nv785_ | new_nv718_ | new_nv818_ | new_nv735_;
  assign new_nv740_ = new_n_n57_ & new_nv732_ & new_nv699_;
  assign new_nv761_ = new_n_n53_ & new_nv699_ & new_nv749_ & new_nv649_;
  assign new_nv772_ = new_n_n59_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv781_ = new_n_n50_ & new_nv699_ & new_nv652_ & new_nv649_ & new_nv706_;
  assign new_nv791_ = new_n_n277_ & new_n_n56_ & new_nv649_ & new_nv627_ & new_nv699_ & new_nv652_;
  assign new_nv802_ = new_nv799_ & new_nv627_ & new_n_n169_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv811_ = new_nv799_ & new_nv627_ & new_n_n160_ & new_nv652_ & new_nv1316_ & new_nv699_ & new_nv649_;
  assign new_nv821_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n210_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv830_ = new_nv1316_ & new_nv652_ & new_nv1315_ & new_nv1310_ & new_nv1287_ & new_n_n280_ & new_nv1263_ & new_nv1316_ & new_n_n281_ & new_n_n201_ & new_nv627_ & new_nv660_ & new_nv649_ & new_nv699_;
  assign new_nv840_ = new_n_n25_ & new_nv831_;
  assign new_nv858_ = new_n_n7_ & new_nv831_;
  assign new_n_n116_ = new_nv935_ | new_nv901_ | new_nv1002_ | new_nv969_ | new_nv833_ | new_nv1035_ | new_nv867_;
  assign new_nv872_ = new_n_n27_ & new_nv865_ & new_nv864_;
  assign new_n_n107_ = new_nv944_ | new_nv910_ | new_nv1011_ | new_nv978_ | new_nv842_ | new_nv1044_ | new_nv876_;
  assign new_nv881_ = new_n_n18_ & new_nv865_ & new_nv864_;
  assign new_n_n98_ = new_nv953_ | new_nv919_ | new_nv1020_ | new_nv987_ | new_nv851_ | new_nv1053_ | new_nv885_;
  assign new_nv890_ = new_n_n9_ & new_nv865_ & new_nv864_;
  assign new_n_n89_ = new_nv962_ | new_nv928_ | new_nv1029_ | new_nv996_ | new_nv860_ | new_nv1062_ | new_nv894_;
  assign new_nv902_ = new_n_n31_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv911_ = new_n_n22_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv929_ = new_n_n4_ & new_nv864_ & new_nv899_ & new_nv898_;
  assign new_nv940_ = new_n_n27_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv949_ = new_n_n18_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv958_ = new_n_n9_ & new_nv864_ & new_nv932_ & new_nv898_ & new_nv933_;
  assign new_nv969_ = new_nv967_ & new_n_n32_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv978_ = new_nv967_ & new_n_n23_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv987_ = new_nv967_ & new_n_n14_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv996_ = new_nv967_ & new_n_n5_ & new_nv898_ & new_nv966_ & new_nv864_ & new_nv932_;
  assign new_nv1006_ = new_n_n277_ & new_nv966_ & new_n_n28_ & new_nv932_ & new_nv1000_ & new_nv864_ & new_nv898_;
  assign new_nv1034_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n171_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1043_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n162_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1052_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n173_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1061_ = new_nv1000_ & new_nv932_ & new_nv1316_ & new_n_n187_ & new_n_n181_ & new_nv966_ & new_nv1316_ & new_nv898_ & new_nv864_;
  assign new_nv1071_ = new_n_n211_ & new_nv1066_;
  assign new_nv1080_ = new_n_n202_ & new_nv1066_;
  assign new_n_n82_ = new_nv1103_ | new_nv1122_ | new_nv1117_ | new_nv1087_ | new_nv1070_;
  assign new_nv1092_ = new_n_n207_ & new_nv1083_ & new_nv1082_;
  assign new_nv556_ = ~new_nv554_;
  assign new_nv1124_ = new_nv1316_ & new_n_n187_ & new_n_n179_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_n_n70_ = new_nv1147_ | new_nv1144_ | new_nv1141_ | new_nv1149_ | new_nv1135_;
  assign new_nv560_ = new_nv1316_ & new_nv1315_ & new_nv1310_;
  assign new_nv749_ = new_nv1315_ & new_nv1287_ & new_n_n282_;
  assign new_nv1139_ = new_nv1316_ & new_n_n281_ & new_n_n280_;
  assign new_nv1123_ = new_nv1316_ & new_n_n187_ & new_n_n177_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1141_ = new_n_n155_ & new_nv1136_ & new_nv1140_ & new_nv660_ & new_n_n277_;
  assign new_nv557_ = new_nv1316_ & new_nv1295_ & new_n_n275_ & new_nv1315_;
  assign new_nv799_ = new_n_n187_ & new_nv1316_;
  assign new_nv1134_ = new_nv1316_ & new_nv1302_ & new_n_n275_ & new_nv1315_;
  assign new_nv1122_ = new_nv1316_ & new_n_n187_ & new_n_n178_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1144_ = new_nv1143_ & new_nv1136_ & new_nv1140_ & new_nv660_ & new_nv1316_;
  assign new_nv573_ = new_nv1315_ & new_nv1302_ & new_n_n275_;
  assign new_nv706_ = new_n_n275_ & new_nv1315_;
  assign new_nv1116_ = new_nv1315_ & new_n_n278_ & new_nv1310_ & new_nv1300_ & new_nv1295_ & new_nv1309_ & new_nv1299_ & new_nv1316_;
  assign new_nv1121_ = new_nv1316_ & new_n_n187_ & new_n_n176_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1147_ = new_nv582_ & new_nv1146_ & new_nv660_ & new_nv1316_ & new_nv1136_ & new_nv1140_;
  assign new_nv569_ = new_nv1315_ & new_n_n280_ & new_n_n281_ & new_nv1302_ & new_nv1287_;
  assign new_nv732_ = new_nv1315_ & new_nv1295_ & new_nv1287_ & new_nv1289_;
  assign new_nv1083_ = new_nv1315_ & new_nv1295_ & new_n_n275_ & new_nv1309_;
  assign new_nv421_ = ~new_n_n68_;
  assign new_nv259_ = new_n_n250_ & new_n_n68_;
  assign new_n_n63_ = new_nv325_ | new_nv553_ | new_nv357_ | new_nv270_ | new_nv237_;
  assign new_nv383_ = new_n_n219_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv1120_ = new_nv1316_ & new_n_n187_ & new_n_n173_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1310_ = ~new_n_n275_;
  assign new_nv1155_ = ~new_nv1153_;
  assign new_nv864_ = ~new_nv831_;
  assign new_nv586_ = ~new_nv1146_;
  assign new_nv260_ = new_n_n249_ & new_n_n68_;
  assign new_nv270_ = new_n_n264_ & new_n_n67_ & new_nv421_;
  assign new_nv373_ = new_n_n229_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv1119_ = new_nv1316_ & new_n_n187_ & new_n_n174_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1309_ = ~new_n_n281_;
  assign new_nv1263_ = ~new_n_n282_;
  assign new_nv699_ = ~new_nv697_;
  assign new_nv590_ = ~new_nv587_;
  assign new_nv239_ = new_n_n270_ & new_n_n68_;
  assign new_nv250_ = new_n_n259_ & new_n_n68_;
  assign new_nv363_ = new_n_n251_ & new_nv421_ & new_nv519_ & new_nv486_ & new_n_n65_;
  assign new_nv1302_ = ~new_n_n274_;
  assign new_nv1140_ = ~new_nv1139_;
  assign new_nv932_ = ~new_nv899_;
  assign new_nv600_ = ~new_nv631_;
  assign new_nv240_ = new_n_n269_ & new_n_n68_;
  assign new_nv249_ = new_n_n260_ & new_n_n68_;
  assign new_nv341_ = new_n_n245_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv1300_ = ~new_n_n150_;
  assign new_nv1152_ = ~new_nv1150_;
  assign new_nv898_ = ~new_nv865_;
  assign new_nv624_ = ~new_nv622_;
  assign new_nv230_ = new_nv1316_ & new_nv1309_ & new_nv1288_ & new_nv1295_ & new_nv1289_;
  assign new_nv331_ = new_n_n255_ & new_nv421_ & new_n_n66_ & new_nv486_;
  assign new_nv587_ = new_nv1316_ & new_nv1295_ & new_nv1310_ & new_nv1315_;
  assign new_nv865_ = new_n_n279_ & new_nv1299_ & new_nv1309_ & new_nv1315_ & new_n_n278_;
  assign new_nv1150_ = new_nv1316_ & new_nv1315_ & new_n_n275_;
  assign new_nv1288_ = ~new_n_n278_;
  assign new_nv1000_ = ~new_nv967_;
  assign new_nv627_ = ~new_nv706_;
  assign new_nv229_ = new_nv1316_ & new_nv1309_ & new_n_n274_ & new_n_n280_;
  assign new_n_n36_ = new_nv264_ | new_nv504_ | new_nv553_ | new_nv384_;
  assign new_nv622_ = new_nv1287_ & new_nv1315_;
  assign new_nv831_ = new_nv1315_ & new_nv1289_ & new_nv1309_ & new_nv1288_ & new_nv1287_;
  assign new_nv1153_ = new_nv1316_ & new_n_n280_ & new_nv1315_ & new_n_n281_;
  assign new_nv1289_ = ~new_n_n276_;
  assign new_nv966_ = ~new_nv933_;
  assign new_nv646_ = ~new_nv644_;
  assign new_nv310_ = new_n_n244_ & new_n_n67_ & new_nv421_;
  assign new_nv1129_ = new_nv1316_ & new_n_n187_ & new_n_n181_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1151_ = new_n_n154_ & new_nv1150_;
  assign new_nv1316_ = ~new_n_n277_;
  assign new_nv1276_ = ~new_n_n279_;
  assign new_nv1099_ = ~new_nv1083_;
  assign new_nv649_ = ~new_nv732_;
  assign new_nv300_ = new_n_n249_ & new_n_n67_ & new_nv421_;
  assign new_nv1130_ = new_nv1316_ & new_n_n187_ & new_n_n180_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1149_ = new_nv582_ & new_nv586_ & new_nv660_ & new_nv1316_ & new_nv1136_ & new_nv1140_;
  assign new_nv1315_ = ~new_n_n187_;
  assign new_nv1287_ = ~new_n_n152_;
  assign new_nv1082_ = ~new_nv1066_;
  assign new_nv652_ = ~new_nv749_;
  assign new_nv290_ = new_n_n254_ & new_n_n67_ & new_nv421_;
  assign new_nv1128_ = new_nv1316_ & new_n_n187_ & new_n_n182_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1131_ = new_nv1316_ & new_n_n187_ & new_n_n188_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_n_n69_ = new_nv1156_ | new_nv1154_ | new_nv1151_;
  assign new_nv694_ = new_nv1315_ & new_nv1295_ & new_nv1287_ & new_nv1309_;
  assign new_nv1066_ = new_nv1288_ & new_nv1315_ & new_nv1295_ & new_nv1309_ & new_nv1289_ & new_nv1287_;
  assign new_nv1136_ = ~new_nv1134_;
  assign new_nv660_ = ~new_nv799_;
  assign new_nv280_ = new_n_n259_ & new_n_n67_ & new_nv421_;
  assign new_nv1127_ = new_nv1316_ & new_n_n187_ & new_n_n183_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1132_ = new_nv1316_ & new_n_n187_ & new_n_n186_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1154_ = new_nv1153_ & new_nv1152_;
  assign new_nv697_ = new_nv1315_ & new_nv1289_ & new_nv1287_ & new_nv1309_;
  assign new_nv967_ = new_nv1315_ & new_nv1309_ & new_n_n275_;
  assign new_nv1118_ = ~new_nv1116_;
  assign new_nv696_ = ~new_nv694_;
  assign new_nv1126_ = new_nv1316_ & new_n_n187_ & new_n_n184_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1133_ = new_nv1316_ & new_n_n187_ & new_n_n192_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv554_ = new_nv1316_ & new_nv1315_ & new_n_n275_ & new_nv1309_;
  assign new_nv631_ = new_nv1315_ & new_nv1289_ & new_nv1287_;
  assign new_nv933_ = new_nv1289_ & new_nv1315_ & new_n_n280_ & new_n_n281_ & new_n_n282_ & new_nv1287_;
  assign new_nv1143_ = new_nv1316_ & new_nv1315_ & new_n_n274_;
  assign new_nv1295_ = ~new_n_n280_;
  assign new_nv1125_ = new_nv1316_ & new_n_n187_ & new_n_n185_ & new_nv1099_ & new_nv1118_ & new_nv1082_ & new_nv1316_;
  assign new_nv1135_ = new_n_n156_ & new_nv1134_;
  assign new_nv1156_ = new_n_n153_ & new_nv1152_ & new_n_n277_ & new_nv1155_;
  assign new_nv644_ = new_nv1315_ & new_nv1309_ & new_nv1287_;
  assign new_nv899_ = new_nv1276_ & new_nv1315_ & new_n_n278_ & new_nv1309_;
  assign new_nv1146_ = new_nv1316_ & new_nv1315_ & new_nv1310_ & new_nv1309_;
  assign new_nv1299_ = ~new_n_n151_;
endmodule


